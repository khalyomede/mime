module mime

pub enum Mime {
    application_vnd_lotus_1_2_3
    text_vnd_in3d_3dml
    video_3gpp2
    image_avif
    image_avif_sequence
    application_x_krita
    image_heic
    video_3gpp
    audio_3gpp2
    application_x_7z_compressed
    application_octet_stream
    application_x_authorware_bin
    image_x_icns
    audio_mp4
    audio_aac
    audio_mp4a_latm
    audio_aacp
    application_x_authorware_map
    application_x_authorware_seg
    application_x_abiword
    application_vnd_americandynamics_acc
    application_x_ace_compressed
    application_vnd_acucobol
    application_vnd_acucorp
    audio_adpcm
    application_vnd_audiograph
    application_x_font_type1
    application_vnd_ibm_modcap
    application_postscript
    application_vnd_adobe_air_application_installer_package_zip
    application_vnd_amiga_ami
    application_vnd_android_package_archive
    application_x_ms_application
    application_vnd_lotus_approach
    application_pgp_signature
    video_x_ms_asf
    text_x_asm
    application_vnd_accpac_simply_aso
    application_atom_xml
    application_atomcat_xml
    application_atomsvc_xml
    application_vnd_antix_game_component
    audio_basic
    video_x_msvideo
    application_applixware
    application_vnd_airzip_filesecure_azf
    application_vnd_airzip_filesecure_azs
    application_vnd_amazon_ebook
    application_x_msdownload
    application_x_bcpio
    application_x_font_bdf
    application_vnd_syncml_dm_wbxml
    application_vnd_fujitsu_oasysprs
    application_vnd_bmi
    image_bmp
    application_vnd_framemaker
    application_vnd_previewsystems_box
    application_x_bzip2
    image_prs_btif
    application_x_bzip
    text_x_c
    application_vnd_clonk_c4group
    application_vnd_ms_cab_compressed
    application_vnd_curl_car
    application_vnd_ms_pki_seccat
    application_x_director
    application_ccxml_xml
    application_vnd_contact_cmsg
    application_x_netcdf
    application_vnd_mediastation_cdkey
    chemical_x_cdx
    application_vnd_chemdraw_xml
    application_vnd_cinderella
    application_pkix_cert
    image_cgm
    application_x_chat
    application_vnd_ms_htmlhelp
    application_vnd_kde_kchart
    chemical_x_cif
    application_vnd_anser_web_certificate_issue_initiation
    application_vnd_ms_artgalry
    application_vnd_claymore
    application_java_vm
    application_vnd_crick_clicker_keyboard
    application_vnd_crick_clicker_palette
    application_vnd_crick_clicker_template
    application_vnd_crick_clicker_wordbank
    application_vnd_crick_clicker
    application_x_msclip
    application_vnd_cosmocaller
    chemical_x_cmdf
    chemical_x_cml
    application_vnd_yellowriver_custom_menu
    image_x_cmx
    application_vnd_rim_cod
    text_plain
    application_vnd_debian_binary_package
    text_markdown
    application_wasm
    application_x_cpio
    application_mac_compactpro
    application_x_mscardfile
    application_pkix_crl
    application_x_x509_ca_cert
    application_x_csh
    chemical_x_csml
    application_vnd_commonspace
    text_css
    text_csv
    application_cu_seeme
    text_vnd_curl
    application_prs_cww
    application_vnd_mobius_daf
    application_vnd_fdsn_seed
    application_davmount_xml
    text_vnd_curl_dcurl
    application_vnd_oma_dd2_xml
    application_vnd_fujixerox_ddd
    application_x_debian_package
    application_vnd_dreamfactory
    application_vnd_mobius_dis
    image_vnd_djvu
    application_vnd_dna
    application_msword
    application_vnd_ms_word_document_macroenabled_12
    application_vnd_openxmlformats_officedocument_wordprocessingml_document
    application_vnd_ms_word_template_macroenabled_12
    application_vnd_openxmlformats_officedocument_wordprocessingml_template
    application_vnd_osgi_dp
    application_vnd_dpgraph
    text_prs_lines_tag
    application_x_dtbook_xml
    application_xml_dtd
    audio_vnd_dts
    audio_vnd_dts_hd
    application_x_dvi
    model_vnd_dwf
    image_vnd_dwg
    image_vnd_dxf
    application_vnd_spotfire_dxp
    audio_vnd_nuera_ecelp4800
    audio_vnd_nuera_ecelp7470
    audio_vnd_nuera_ecelp9600
    application_ecmascript
    application_vnd_novadigm_edm
    application_vnd_novadigm_edx
    application_vnd_picsel
    application_vnd_pg_osasli
    message_rfc822
    application_emma_xml
    audio_vnd_digital_winds
    application_vnd_ms_fontobject
    application_epub_zip
    application_vnd_eszigno3_xml
    application_vnd_epson_esf
    text_x_setext
    application_vnd_novadigm_ext
    application_andrew_inset
    application_vnd_ezpix_album
    application_vnd_ezpix_package
    text_x_fortran
    video_x_f4v
    image_vnd_fastbidsheet
    application_vnd_fdf
    application_vnd_denovo_fcselayout_link
    application_vnd_fujitsu_oasysgp
    image_x_freehand
    application_x_xfig
    video_x_fli
    application_vnd_micrografx_flo
    video_x_flv
    application_vnd_kde_kivio
    text_vnd_fmi_flexstor
    text_vnd_fly
    application_vnd_frogans_fnc
    image_vnd_fpx
    application_vnd_fsc_weblaunch
    image_vnd_fst
    application_vnd_fluxtime_clip
    application_vnd_anser_web_funds_transfer_initiation
    video_vnd_fvt
    application_vnd_fuzzysheet
    image_g3fax
    application_vnd_groove_account
    model_vnd_gdl
    application_vnd_dynageo
    application_vnd_geometry_explorer
    application_vnd_geogebra_file
    application_vnd_geogebra_tool
    application_vnd_groove_help
    image_gif
    application_vnd_groove_identity_message
    application_vnd_gmx
    application_x_gnumeric
    application_vnd_flographit
    application_vnd_grafeq
    application_srgs
    application_vnd_groove_injector
    application_srgs_xml
    application_x_font_ghostscript
    application_x_gtar
    application_vnd_groove_tool_message
    model_vnd_gtw
    text_vnd_graphviz
    application_x_gzip
    application_gzip
    video_h261
    gcode
    video_h263
    video_h264
    application_vnd_hbci
    application_vnd_gerber
    application_x_hdf
    application_winhlp
    application_vnd_hp_hpgl
    application_vnd_hp_hpid
    application_vnd_hp_hps
    application_mac_binhex40
    application_vnd_kenameaapp
    text_html
    application_vnd_yamaha_hv_dic
    application_vnd_yamaha_hv_voice
    application_vnd_yamaha_hv_script
    application_vnd_iccprofile
    x_conference_x_cooltalk
    image_x_icon
    text_calendar
    image_ief
    application_vnd_shana_informed_formdata
    model_iges
    application_vnd_igloader
    application_vnd_micrografx_igx
    application_vnd_shana_informed_interchange
    application_vnd_accpac_simply_imp
    application_vnd_ms_ims
    application_vnd_shana_informed_package
    application_vnd_ibm_rights_management
    application_vnd_irepository_package_xml
    application_vnd_shana_informed_formtemplate
    application_vnd_immervision_ivp
    application_vnd_immervision_ivu
    text_vnd_sun_j2me_app_descriptor
    application_vnd_jam
    application_java_archive
    text_x_java_source
    application_vnd_jisp
    application_vnd_hp_jlyt
    application_x_java_jnlp_file
    application_vnd_joost_joda_archive
    image_jpeg
    image_pjpeg
    video_jpm
    video_jpeg
    application_x_trash
    application_x_shellscript
    text_javascript
    application_json
    audio_midi
    audio_aiff
    audio_opus
    application_vnd_kde_karbon
    application_vnd_kde_kformula
    application_vnd_kidspiration
    application_x_killustrator
    application_vnd_google_earth_kml_xml
    application_vnd_google_earth_kmz
    application_vnd_kinar
    application_vnd_kde_kontour
    application_vnd_kde_kpresenter
    application_vnd_kde_kspread
    application_vnd_kahootz
    application_vnd_kde_kword
    application_x_latex
    application_vnd_llamagraphics_life_balance_desktop
    application_vnd_llamagraphics_life_balance_exchange_xml
    application_vnd_hhe_lesson_player
    application_vnd_route66_link66_xml
    application_lost_xml
    application_vnd_ms_lrm
    application_vnd_frogans_ltf
    audio_vnd_lucent_voice
    application_vnd_lotus_wordpro
    application_x_msmediaview
    video_mpeg
    audio_mpeg
    audio_x_mpegurl
    video_vnd_mpegurl
    video_x_m4v
    application_mathematica
    application_vnd_ecowin_chart
    text_troff
    application_mathml_xml
    text_mathml
    application_vnd_sqlite3
    application_vnd_mobius_mbk
    application_mbox
    application_vnd_medcalcdata
    application_vnd_mcd
    text_vnd_curl_mcurl
    application_x_msaccess
    image_vnd_ms_modi
    model_mesh
    application_vnd_mfmp
    application_vnd_proteus_magazine
    application_vnd_mif
    video_mj2
    application_vnd_dolby_mlp
    application_vnd_chipnuts_karaoke_mmd
    application_vnd_smaf
    image_vnd_fujixerox_edmics_mmr
    application_x_msmoney
    application_x_mobipocket_ebook
    video_quicktime
    video_x_sgi_movie
    video_mp4
    application_x_iso9660_image
    application_yaml
    application_mp4
    application_vnd_mophun_certificate
    application_vnd_apple_installer_xml
    application_vnd_blueice_multipass
    application_vnd_mophun_application
    application_vnd_ms_project
    application_vnd_ibm_minipay
    application_vnd_mobius_mqy
    application_marc
    application_mediaservercontrol_xml
    application_vnd_fdsn_mseed
    application_vnd_mseq
    application_vnd_epson_msf
    application_vnd_mobius_msl
    application_vnd_muvee_style
    model_vnd_mts
    application_vnd_musician
    application_vnd_recordare_musicxml_xml
    application_vnd_mfer
    application_mxf
    application_vnd_recordare_musicxml
    application_xv_xml
    application_vnd_triscape_mxs
    application_vnd_nokia_n_gage_symbian_install
    application_x_dtbncx_xml
    application_vnd_nokia_n_gage_data
    application_vnd_neurolanguage_nlu
    application_vnd_enliven
    application_vnd_noblenet_directory
    application_vnd_noblenet_sealer
    application_vnd_noblenet_web
    image_vnd_net_fpx
    application_vnd_lotus_notes
    application_vnd_fujitsu_oasys2
    application_vnd_fujitsu_oasys3
    application_vnd_fujitsu_oasys
    application_x_msbinder
    application_oda
    application_vnd_oasis_opendocument_database
    application_vnd_oasis_opendocument_chart
    application_vnd_oasis_opendocument_formula
    application_vnd_oasis_opendocument_formula_template
    application_vnd_oasis_opendocument_graphics
    application_vnd_oasis_opendocument_image
    application_vnd_oasis_opendocument_presentation
    application_vnd_oasis_opendocument_spreadsheet
    application_vnd_oasis_opendocument_text
    audio_ogg
    video_x_matroska
    audio_x_matroska
    video_ogg
    application_ogg
    application_onenote
    application_oebps_package_xml
    application_vnd_palm
    application_vnd_lotus_organizer
    application_vnd_yamaha_openscoreformat
    application_vnd_yamaha_openscoreformat_osfpvg_xml
    application_vnd_oasis_opendocument_chart_template
    font_woff
    font_woff2
    application_x_redhat_package_manager
    application_x_perl
    audio_webm
    video_webm
    image_webp
    application_x_font_otf
    font_otf
    application_vnd_oasis_opendocument_graphics_template
    application_vnd_oasis_opendocument_text_web
    application_vnd_oasis_opendocument_image_template
    application_vnd_oasis_opendocument_text_master
    application_vnd_oasis_opendocument_presentation_template
    application_vnd_oasis_opendocument_spreadsheet_template
    application_vnd_oasis_opendocument_text_template
    application_vnd_openofficeorg_extension
    text_x_pascal
    application_pkcs10
    application_x_pkcs12
    application_x_pkcs7_certificates
    application_pkcs7_mime
    application_x_pkcs7_certreqresp
    application_pkcs7_signature
    application_vnd_powerbuilder6
    image_x_portable_bitmap
    application_x_font_pcf
    application_vnd_hp_pcl
    application_vnd_hp_pclxl
    image_x_pict
    application_vnd_curl_pcurl
    image_x_pcx
    application_pdf
    application_font_tdpfr
    image_x_portable_graymap
    application_x_chess_pgn
    application_pgp_encrypted
    application_pkixcmp
    application_pkix_pkipath
    application_vnd_3gpp_pic_bw_large
    application_vnd_mobius_plc
    application_vnd_pocketlearn
    application_pls_xml
    application_vnd_ctc_posml
    image_png
    image_x_portable_anymap
    application_vnd_macports_portpkg
    application_vnd_ms_powerpoint
    application_vnd_ms_powerpoint_template_macroenabled_12
    application_vnd_openxmlformats_officedocument_presentationml_template
    application_vnd_ms_powerpoint_addin_macroenabled_12
    application_vnd_cups_ppd
    image_x_portable_pixmap
    application_vnd_ms_powerpoint_slideshow_macroenabled_12
    application_vnd_openxmlformats_officedocument_presentationml_slideshow
    application_vnd_ms_powerpoint_presentation_macroenabled_12
    application_vnd_openxmlformats_officedocument_presentationml_presentation
    application_vnd_lotus_freelance
    application_pics_rules
    application_prql
    application_vnd_3gpp_pic_bw_small
    image_vnd_adobe_photoshop
    application_x_font_linux_psf
    application_vnd_pvi_ptid1
    application_x_mspublisher
    application_vnd_3gpp_pic_bw_var
    application_vnd_3m_post_it_notes
    text_x_python
    audio_vnd_ms_playready_media_pya
    video_vnd_ms_playready_media_pyv
    application_vnd_epson_quickanime
    application_vnd_intu_qbo
    application_vnd_intu_qfx
    application_vnd_publishare_delta_tree
    application_vnd_quark_quarkxpress
    audio_x_pn_realaudio
    application_vnd_rar
    application_x_rar_compressed
    image_x_cmu_raster
    application_vnd_ipunplugged_rcprofile
    application_rdf_xml
    application_vnd_data_vision_rdz
    application_vnd_businessobjects
    application_x_dtbresource_xml
    image_x_rgb
    application_reginfo_xml
    application_resource_lists_xml
    image_vnd_fujixerox_edmics_rlc
    application_resource_lists_diff_xml
    application_vnd_rn_realmedia
    audio_x_pn_realaudio_plugin
    application_vnd_jcp_javame_midlet_rms
    application_relax_ng_compact_syntax
    application_x_rpm
    application_vnd_nokia_radio_presets
    application_vnd_nokia_radio_preset
    application_sparql_query
    application_rls_services_xml
    application_rsd_xml
    application_rss_xml
    application_rtf
    text_richtext
    application_vnd_yamaha_smaf_audio
    application_sbml_xml
    application_vnd_ibm_secure_container
    application_x_msschedule
    application_vnd_lotus_screencam
    application_scvp_cv_request
    application_scvp_cv_response
    text_vnd_curl_scurl
    application_vnd_stardivision_draw
    application_vnd_stardivision_calc
    application_vnd_stardivision_impress
    application_vnd_solent_sdkm_xml
    application_sdp
    application_vnd_stardivision_writer
    application_vnd_seemail
    application_vnd_sema
    application_vnd_semd
    application_vnd_semf
    application_java_serialized_object
    application_set_payment_initiation
    application_set_registration_initiation
    application_vnd_hydrostatix_sof_data
    application_vnd_spotfire_sfs
    application_vnd_stardivision_writer_global
    text_sgml
    application_x_sh
    application_x_shar
    application_shf_xml
    text_vnd_wap_si
    application_vnd_wap_sic
    application_vnd_symbian_install
    application_x_stuffit
    application_x_stuffitx
    application_vnd_koan
    text_vnd_wap_sl
    application_vnd_wap_slc
    application_vnd_ms_powerpoint_slide_macroenabled_12
    application_vnd_openxmlformats_officedocument_presentationml_slide
    application_vnd_epson_salt
    application_vnd_stardivision_math
    application_smil_xml
    application_x_font_snf
    application_vnd_yamaha_smaf_phrase
    application_x_futuresplash
    text_vnd_in3d_spot
    application_scvp_vp_response
    application_scvp_vp_request
    application_x_wais_source
    application_sparql_results_xml
    application_vnd_kodak_descriptor
    application_vnd_epson_ssf
    application_ssml_xml
    application_vnd_sun_xml_calc_template
    application_vnd_sun_xml_draw_template
    application_vnd_wt_stf
    application_vnd_sun_xml_impress_template
    application_hyperstudio
    application_vnd_ms_pki_stl
    application_vnd_pg_format
    application_vnd_sun_xml_writer_template
    application_vnd_sus_calendar
    application_x_sv4cpio
    application_x_sv4crc
    application_vnd_svd
    image_svg_xml
    application_x_shockwave_flash
    application_vnd_arastra_swi
    application_vnd_sun_xml_calc
    application_vnd_sun_xml_draw
    application_vnd_sun_xml_writer_global
    application_vnd_sun_xml_impress
    application_vnd_sun_xml_math
    application_vnd_sun_xml_writer
    application_vnd_tao_intent_module_archive
    application_x_tar
    application_vnd_3gpp2_tcap
    application_x_tcl
    application_vnd_smart_teacher
    application_x_tex
    application_x_texinfo
    application_x_tex_tfm
    image_tiff
    application_vnd_tmobile_livetv
    application_x_bittorrent
    application_vnd_groove_tool_template
    application_vnd_trid_tpt
    application_vnd_trueapp
    application_x_msterminal
    text_tab_separated_values
    application_x_font_ttf
    application_vnd_simtech_mindmapper
    application_vnd_genomatix_tuxedo
    application_vnd_mobius_txf
    application_vnd_ufdl
    test_mimetype
    application_vnd_umajin
    application_vnd_unity
    application_vnd_uoml_xml
    text_uri_list
    application_x_ustar
    application_vnd_uiq_theme
    text_x_uuencode
    application_x_cdlink
    text_x_vcard
    application_vnd_groove_vcard
    text_x_vcalendar
    application_vnd_vcx
    application_vnd_visionary
    video_vnd_vivo
    model_vrml
    application_vnd_visio
    application_vnd_vsf
    model_vnd_vtu
    application_voicexml_xml
    application_x_doom
    video_mp2t
    audio_vnd_wav
    audio_x_ms_wax
    image_vnd_wap_wbmp
    application_vnd_criticaltools_wbs_xml
    application_vnd_wap_wbxml
    application_vnd_ms_works
    video_x_ms_wm
    audio_x_ms_wma
    application_x_ms_wmd
    application_x_msmetafile
    text_vnd_wap_wml
    application_vnd_wap_wmlc
    text_vnd_wap_wmlscript
    application_vnd_wap_wmlscriptc
    video_x_ms_wmv
    video_x_ms_wmx
    application_x_ms_wmz
    application_vnd_wordperfect
    application_vnd_ms_wpl
    application_vnd_wqd
    application_x_mswrite
    application_wsdl_xml
    application_wspolicy_xml
    application_vnd_webturbo
    video_x_ms_wvx
    application_vnd_hzn_3d_crossword
    application_x_silverlight_app
    application_vnd_xara
    application_x_ms_xbap
    application_vnd_fujixerox_docuworks_binder
    image_x_xbitmap
    application_vnd_syncml_dm_xml
    application_vnd_adobe_xdp_xml
    application_vnd_fujixerox_docuworks
    application_xenc_xml
    application_patch_ops_error_xml
    application_vnd_adobe_xfdf
    application_vnd_xfdl
    application_xhtml_xml
    image_vnd_xiff
    application_vnd_ms_excel
    application_vnd_ms_excel_addin_macroenabled_12
    application_vnd_ms_excel_sheet_binary_macroenabled_12
    application_vnd_ms_excel_sheet_macroenabled_12
    application_vnd_openxmlformats_officedocument_spreadsheetml_sheet
    application_vnd_ms_excel_template_macroenabled_12
    application_vnd_openxmlformats_officedocument_spreadsheetml_template
    application_xml
    application_vnd_olpc_sugar
    application_xop_xml
    application_x_xpinstall
    image_x_xpixmap
    application_vnd_is_xpr
    application_vnd_ms_xpsdocument
    application_vnd_intercon_formnet
    application_xslt_xml
    application_vnd_syncml_xml
    application_xspf_xml
    application_vnd_mozilla_xul_xml
    image_x_xwindowdump
    chemical_x_xyz
    application_vnd_zzazz_deck_xml
    application_zip
    application_x_zip_compressed
    application_zip_compressed
    application_vnd_zul
    application_vnd_handheld_entertainment_xml
    image_x_adobe_dng
    image_x_sony_arw
    image_x_canon_cr2
    image_x_canon_crw
    image_x_kodak_dcr
    image_x_epson_erf
    image_x_kodak_k25
    image_x_kodak_kdc
    image_x_minolta_mrw
    image_x_nikon_nef
    image_x_olympus_orf
    image_x_pentax_pef
    image_x_fuji_raf
    image_x_panasonic_raw
    audio_flac
    image_x_sony_sr2
    image_x_sony_srf
    image_x_sigma_x3f
}
