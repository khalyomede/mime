module mime

pub fn Mime.from_text(text string) ?Mime {
    return match text {
        'application/vnd.lotus-1-2-3' { Mime.application_vnd_lotus_1_2_3 }
        'text/vnd.in3d.3dml' { Mime.text_vnd_in3d_3dml }
        'video/3gpp2' { Mime.video_3gpp2 }
        'image/avif' { Mime.image_avif }
        'image/avif-sequence' { Mime.image_avif_sequence }
        'application/x-krita' { Mime.application_x_krita }
        'image/heic' { Mime.image_heic }
        'video/3gpp' { Mime.video_3gpp }
        'audio/3gpp2' { Mime.audio_3gpp2 }
        'application/x-7z-compressed' { Mime.application_x_7z_compressed }
        'application/octet-stream' { Mime.application_octet_stream }
        'application/x-authorware-bin' { Mime.application_x_authorware_bin }
        'image/x-icns' { Mime.image_x_icns }
        'audio/mp4' { Mime.audio_mp4 }
        'audio/aac' { Mime.audio_aac }
        'audio/mp4a-latm' { Mime.audio_mp4a_latm }
        'audio/aacp' { Mime.audio_aacp }
        'application/x-authorware-map' { Mime.application_x_authorware_map }
        'application/x-authorware-seg' { Mime.application_x_authorware_seg }
        'application/x-abiword' { Mime.application_x_abiword }
        'application/vnd.americandynamics.acc' { Mime.application_vnd_americandynamics_acc }
        'application/x-ace-compressed' { Mime.application_x_ace_compressed }
        'application/vnd.acucobol' { Mime.application_vnd_acucobol }
        'application/vnd.acucorp' { Mime.application_vnd_acucorp }
        'audio/adpcm' { Mime.audio_adpcm }
        'application/vnd.audiograph' { Mime.application_vnd_audiograph }
        'application/x-font-type1' { Mime.application_x_font_type1 }
        'application/vnd.ibm.modcap' { Mime.application_vnd_ibm_modcap }
        'application/postscript' { Mime.application_postscript }
        'application/vnd.adobe.air-application-installer-package+zip' { Mime.application_vnd_adobe_air_application_installer_package_zip }
        'application/vnd.amiga.ami' { Mime.application_vnd_amiga_ami }
        'application/vnd.android.package-archive' { Mime.application_vnd_android_package_archive }
        'application/x-ms-application' { Mime.application_x_ms_application }
        'application/vnd.lotus-approach' { Mime.application_vnd_lotus_approach }
        'application/pgp-signature' { Mime.application_pgp_signature }
        'video/x-ms-asf' { Mime.video_x_ms_asf }
        'text/x-asm' { Mime.text_x_asm }
        'application/vnd.accpac.simply.aso' { Mime.application_vnd_accpac_simply_aso }
        'application/atom+xml' { Mime.application_atom_xml }
        'application/atomcat+xml' { Mime.application_atomcat_xml }
        'application/atomsvc+xml' { Mime.application_atomsvc_xml }
        'application/vnd.antix.game-component' { Mime.application_vnd_antix_game_component }
        'audio/basic' { Mime.audio_basic }
        'video/x-msvideo' { Mime.video_x_msvideo }
        'application/applixware' { Mime.application_applixware }
        'application/vnd.airzip.filesecure.azf' { Mime.application_vnd_airzip_filesecure_azf }
        'application/vnd.airzip.filesecure.azs' { Mime.application_vnd_airzip_filesecure_azs }
        'application/vnd.amazon.ebook' { Mime.application_vnd_amazon_ebook }
        'application/x-msdownload' { Mime.application_x_msdownload }
        'application/x-bcpio' { Mime.application_x_bcpio }
        'application/x-font-bdf' { Mime.application_x_font_bdf }
        'application/vnd.syncml.dm+wbxml' { Mime.application_vnd_syncml_dm_wbxml }
        'application/vnd.fujitsu.oasysprs' { Mime.application_vnd_fujitsu_oasysprs }
        'application/vnd.bmi' { Mime.application_vnd_bmi }
        'image/bmp' { Mime.image_bmp }
        'application/vnd.framemaker' { Mime.application_vnd_framemaker }
        'application/vnd.previewsystems.box' { Mime.application_vnd_previewsystems_box }
        'application/x-bzip2' { Mime.application_x_bzip2 }
        'image/prs.btif' { Mime.image_prs_btif }
        'application/x-bzip' { Mime.application_x_bzip }
        'text/x-c' { Mime.text_x_c }
        'application/vnd.clonk.c4group' { Mime.application_vnd_clonk_c4group }
        'application/vnd.ms-cab-compressed' { Mime.application_vnd_ms_cab_compressed }
        'application/vnd.curl.car' { Mime.application_vnd_curl_car }
        'application/vnd.ms-pki.seccat' { Mime.application_vnd_ms_pki_seccat }
        'application/x-director' { Mime.application_x_director }
        'application/ccxml+xml' { Mime.application_ccxml_xml }
        'application/vnd.contact.cmsg' { Mime.application_vnd_contact_cmsg }
        'application/x-netcdf' { Mime.application_x_netcdf }
        'application/vnd.mediastation.cdkey' { Mime.application_vnd_mediastation_cdkey }
        'chemical/x-cdx' { Mime.chemical_x_cdx }
        'application/vnd.chemdraw+xml' { Mime.application_vnd_chemdraw_xml }
        'application/vnd.cinderella' { Mime.application_vnd_cinderella }
        'application/pkix-cert' { Mime.application_pkix_cert }
        'image/cgm' { Mime.image_cgm }
        'application/x-chat' { Mime.application_x_chat }
        'application/vnd.ms-htmlhelp' { Mime.application_vnd_ms_htmlhelp }
        'application/vnd.kde.kchart' { Mime.application_vnd_kde_kchart }
        'chemical/x-cif' { Mime.chemical_x_cif }
        'application/vnd.anser-web-certificate-issue-initiation' { Mime.application_vnd_anser_web_certificate_issue_initiation }
        'application/vnd.ms-artgalry' { Mime.application_vnd_ms_artgalry }
        'application/vnd.claymore' { Mime.application_vnd_claymore }
        'application/java-vm' { Mime.application_java_vm }
        'application/vnd.crick.clicker.keyboard' { Mime.application_vnd_crick_clicker_keyboard }
        'application/vnd.crick.clicker.palette' { Mime.application_vnd_crick_clicker_palette }
        'application/vnd.crick.clicker.template' { Mime.application_vnd_crick_clicker_template }
        'application/vnd.crick.clicker.wordbank' { Mime.application_vnd_crick_clicker_wordbank }
        'application/vnd.crick.clicker' { Mime.application_vnd_crick_clicker }
        'application/x-msclip' { Mime.application_x_msclip }
        'application/vnd.cosmocaller' { Mime.application_vnd_cosmocaller }
        'chemical/x-cmdf' { Mime.chemical_x_cmdf }
        'chemical/x-cml' { Mime.chemical_x_cml }
        'application/vnd.yellowriver-custom-menu' { Mime.application_vnd_yellowriver_custom_menu }
        'image/x-cmx' { Mime.image_x_cmx }
        'application/vnd.rim.cod' { Mime.application_vnd_rim_cod }
        'text/plain' { Mime.text_plain }
        'application/vnd.debian.binary-package' { Mime.application_vnd_debian_binary_package }
        'text/markdown' { Mime.text_markdown }
        'application/wasm' { Mime.application_wasm }
        'application/x-cpio' { Mime.application_x_cpio }
        'application/mac-compactpro' { Mime.application_mac_compactpro }
        'application/x-mscardfile' { Mime.application_x_mscardfile }
        'application/pkix-crl' { Mime.application_pkix_crl }
        'application/x-x509-ca-cert' { Mime.application_x_x509_ca_cert }
        'application/x-csh' { Mime.application_x_csh }
        'chemical/x-csml' { Mime.chemical_x_csml }
        'application/vnd.commonspace' { Mime.application_vnd_commonspace }
        'text/css' { Mime.text_css }
        'text/csv' { Mime.text_csv }
        'application/cu-seeme' { Mime.application_cu_seeme }
        'text/vnd.curl' { Mime.text_vnd_curl }
        'application/prs.cww' { Mime.application_prs_cww }
        'application/vnd.mobius.daf' { Mime.application_vnd_mobius_daf }
        'application/vnd.fdsn.seed' { Mime.application_vnd_fdsn_seed }
        'application/davmount+xml' { Mime.application_davmount_xml }
        'text/vnd.curl.dcurl' { Mime.text_vnd_curl_dcurl }
        'application/vnd.oma.dd2+xml' { Mime.application_vnd_oma_dd2_xml }
        'application/vnd.fujixerox.ddd' { Mime.application_vnd_fujixerox_ddd }
        'application/x-debian-package' { Mime.application_x_debian_package }
        'application/vnd.dreamfactory' { Mime.application_vnd_dreamfactory }
        'application/vnd.mobius.dis' { Mime.application_vnd_mobius_dis }
        'image/vnd.djvu' { Mime.image_vnd_djvu }
        'application/vnd.dna' { Mime.application_vnd_dna }
        'application/msword' { Mime.application_msword }
        'application/vnd.ms-word.document.macroenabled.12' { Mime.application_vnd_ms_word_document_macroenabled_12 }
        'application/vnd.openxmlformats-officedocument.wordprocessingml.document' { Mime.application_vnd_openxmlformats_officedocument_wordprocessingml_document }
        'application/vnd.ms-word.template.macroenabled.12' { Mime.application_vnd_ms_word_template_macroenabled_12 }
        'application/vnd.openxmlformats-officedocument.wordprocessingml.template' { Mime.application_vnd_openxmlformats_officedocument_wordprocessingml_template }
        'application/vnd.osgi.dp' { Mime.application_vnd_osgi_dp }
        'application/vnd.dpgraph' { Mime.application_vnd_dpgraph }
        'text/prs.lines.tag' { Mime.text_prs_lines_tag }
        'application/x-dtbook+xml' { Mime.application_x_dtbook_xml }
        'application/xml-dtd' { Mime.application_xml_dtd }
        'audio/vnd.dts' { Mime.audio_vnd_dts }
        'audio/vnd.dts.hd' { Mime.audio_vnd_dts_hd }
        'application/x-dvi' { Mime.application_x_dvi }
        'model/vnd.dwf' { Mime.model_vnd_dwf }
        'image/vnd.dwg' { Mime.image_vnd_dwg }
        'image/vnd.dxf' { Mime.image_vnd_dxf }
        'application/vnd.spotfire.dxp' { Mime.application_vnd_spotfire_dxp }
        'audio/vnd.nuera.ecelp4800' { Mime.audio_vnd_nuera_ecelp4800 }
        'audio/vnd.nuera.ecelp7470' { Mime.audio_vnd_nuera_ecelp7470 }
        'audio/vnd.nuera.ecelp9600' { Mime.audio_vnd_nuera_ecelp9600 }
        'application/ecmascript' { Mime.application_ecmascript }
        'application/vnd.novadigm.edm' { Mime.application_vnd_novadigm_edm }
        'application/vnd.novadigm.edx' { Mime.application_vnd_novadigm_edx }
        'application/vnd.picsel' { Mime.application_vnd_picsel }
        'application/vnd.pg.osasli' { Mime.application_vnd_pg_osasli }
        'message/rfc822' { Mime.message_rfc822 }
        'application/emma+xml' { Mime.application_emma_xml }
        'audio/vnd.digital-winds' { Mime.audio_vnd_digital_winds }
        'application/vnd.ms-fontobject' { Mime.application_vnd_ms_fontobject }
        'application/epub+zip' { Mime.application_epub_zip }
        'application/vnd.eszigno3+xml' { Mime.application_vnd_eszigno3_xml }
        'application/vnd.epson.esf' { Mime.application_vnd_epson_esf }
        'text/x-setext' { Mime.text_x_setext }
        'application/vnd.novadigm.ext' { Mime.application_vnd_novadigm_ext }
        'application/andrew-inset' { Mime.application_andrew_inset }
        'application/vnd.ezpix-album' { Mime.application_vnd_ezpix_album }
        'application/vnd.ezpix-package' { Mime.application_vnd_ezpix_package }
        'text/x-fortran' { Mime.text_x_fortran }
        'video/x-f4v' { Mime.video_x_f4v }
        'image/vnd.fastbidsheet' { Mime.image_vnd_fastbidsheet }
        'application/vnd.fdf' { Mime.application_vnd_fdf }
        'application/vnd.denovo.fcselayout-link' { Mime.application_vnd_denovo_fcselayout_link }
        'application/vnd.fujitsu.oasysgp' { Mime.application_vnd_fujitsu_oasysgp }
        'image/x-freehand' { Mime.image_x_freehand }
        'application/x-xfig' { Mime.application_x_xfig }
        'video/x-fli' { Mime.video_x_fli }
        'application/vnd.micrografx.flo' { Mime.application_vnd_micrografx_flo }
        'video/x-flv' { Mime.video_x_flv }
        'application/vnd.kde.kivio' { Mime.application_vnd_kde_kivio }
        'text/vnd.fmi.flexstor' { Mime.text_vnd_fmi_flexstor }
        'text/vnd.fly' { Mime.text_vnd_fly }
        'application/vnd.frogans.fnc' { Mime.application_vnd_frogans_fnc }
        'image/vnd.fpx' { Mime.image_vnd_fpx }
        'application/vnd.fsc.weblaunch' { Mime.application_vnd_fsc_weblaunch }
        'image/vnd.fst' { Mime.image_vnd_fst }
        'application/vnd.fluxtime.clip' { Mime.application_vnd_fluxtime_clip }
        'application/vnd.anser-web-funds-transfer-initiation' { Mime.application_vnd_anser_web_funds_transfer_initiation }
        'video/vnd.fvt' { Mime.video_vnd_fvt }
        'application/vnd.fuzzysheet' { Mime.application_vnd_fuzzysheet }
        'image/g3fax' { Mime.image_g3fax }
        'application/vnd.groove-account' { Mime.application_vnd_groove_account }
        'model/vnd.gdl' { Mime.model_vnd_gdl }
        'application/vnd.dynageo' { Mime.application_vnd_dynageo }
        'application/vnd.geometry-explorer' { Mime.application_vnd_geometry_explorer }
        'application/vnd.geogebra.file' { Mime.application_vnd_geogebra_file }
        'application/vnd.geogebra.tool' { Mime.application_vnd_geogebra_tool }
        'application/vnd.groove-help' { Mime.application_vnd_groove_help }
        'image/gif' { Mime.image_gif }
        'application/vnd.groove-identity-message' { Mime.application_vnd_groove_identity_message }
        'application/vnd.gmx' { Mime.application_vnd_gmx }
        'application/x-gnumeric' { Mime.application_x_gnumeric }
        'application/vnd.flographit' { Mime.application_vnd_flographit }
        'application/vnd.grafeq' { Mime.application_vnd_grafeq }
        'application/srgs' { Mime.application_srgs }
        'application/vnd.groove-injector' { Mime.application_vnd_groove_injector }
        'application/srgs+xml' { Mime.application_srgs_xml }
        'application/x-font-ghostscript' { Mime.application_x_font_ghostscript }
        'application/x-gtar' { Mime.application_x_gtar }
        'application/vnd.groove-tool-message' { Mime.application_vnd_groove_tool_message }
        'model/vnd.gtw' { Mime.model_vnd_gtw }
        'text/vnd.graphviz' { Mime.text_vnd_graphviz }
        'application/x-gzip' { Mime.application_x_gzip }
        'application/gzip' { Mime.application_gzip }
        'video/h261' { Mime.video_h261 }
        'gcode' { Mime.gcode }
        'video/h263' { Mime.video_h263 }
        'video/h264' { Mime.video_h264 }
        'application/vnd.hbci' { Mime.application_vnd_hbci }
        'application/vnd.gerber' { Mime.application_vnd_gerber }
        'application/x-hdf' { Mime.application_x_hdf }
        'application/winhlp' { Mime.application_winhlp }
        'application/vnd.hp-hpgl' { Mime.application_vnd_hp_hpgl }
        'application/vnd.hp-hpid' { Mime.application_vnd_hp_hpid }
        'application/vnd.hp-hps' { Mime.application_vnd_hp_hps }
        'application/mac-binhex40' { Mime.application_mac_binhex40 }
        'application/vnd.kenameaapp' { Mime.application_vnd_kenameaapp }
        'text/html' { Mime.text_html }
        'application/vnd.yamaha.hv-dic' { Mime.application_vnd_yamaha_hv_dic }
        'application/vnd.yamaha.hv-voice' { Mime.application_vnd_yamaha_hv_voice }
        'application/vnd.yamaha.hv-script' { Mime.application_vnd_yamaha_hv_script }
        'application/vnd.iccprofile' { Mime.application_vnd_iccprofile }
        'x-conference/x-cooltalk' { Mime.x_conference_x_cooltalk }
        'image/x-icon' { Mime.image_x_icon }
        'text/calendar' { Mime.text_calendar }
        'image/ief' { Mime.image_ief }
        'application/vnd.shana.informed.formdata' { Mime.application_vnd_shana_informed_formdata }
        'model/iges' { Mime.model_iges }
        'application/vnd.igloader' { Mime.application_vnd_igloader }
        'application/vnd.micrografx.igx' { Mime.application_vnd_micrografx_igx }
        'application/vnd.shana.informed.interchange' { Mime.application_vnd_shana_informed_interchange }
        'application/vnd.accpac.simply.imp' { Mime.application_vnd_accpac_simply_imp }
        'application/vnd.ms-ims' { Mime.application_vnd_ms_ims }
        'application/vnd.shana.informed.package' { Mime.application_vnd_shana_informed_package }
        'application/vnd.ibm.rights-management' { Mime.application_vnd_ibm_rights_management }
        'application/vnd.irepository.package+xml' { Mime.application_vnd_irepository_package_xml }
        'application/vnd.shana.informed.formtemplate' { Mime.application_vnd_shana_informed_formtemplate }
        'application/vnd.immervision-ivp' { Mime.application_vnd_immervision_ivp }
        'application/vnd.immervision-ivu' { Mime.application_vnd_immervision_ivu }
        'text/vnd.sun.j2me.app-descriptor' { Mime.text_vnd_sun_j2me_app_descriptor }
        'application/vnd.jam' { Mime.application_vnd_jam }
        'application/java-archive' { Mime.application_java_archive }
        'text/x-java-source' { Mime.text_x_java_source }
        'application/vnd.jisp' { Mime.application_vnd_jisp }
        'application/vnd.hp-jlyt' { Mime.application_vnd_hp_jlyt }
        'application/x-java-jnlp-file' { Mime.application_x_java_jnlp_file }
        'application/vnd.joost.joda-archive' { Mime.application_vnd_joost_joda_archive }
        'image/jpeg' { Mime.image_jpeg }
        'image/pjpeg' { Mime.image_pjpeg }
        'video/jpm' { Mime.video_jpm }
        'video/jpeg' { Mime.video_jpeg }
        'application/x-trash' { Mime.application_x_trash }
        'application/x-shellscript' { Mime.application_x_shellscript }
        'text/javascript' { Mime.text_javascript }
        'application/json' { Mime.application_json }
        'audio/midi' { Mime.audio_midi }
        'audio/aiff' { Mime.audio_aiff }
        'audio/opus' { Mime.audio_opus }
        'application/vnd.kde.karbon' { Mime.application_vnd_kde_karbon }
        'application/vnd.kde.kformula' { Mime.application_vnd_kde_kformula }
        'application/vnd.kidspiration' { Mime.application_vnd_kidspiration }
        'application/x-killustrator' { Mime.application_x_killustrator }
        'application/vnd.google-earth.kml+xml' { Mime.application_vnd_google_earth_kml_xml }
        'application/vnd.google-earth.kmz' { Mime.application_vnd_google_earth_kmz }
        'application/vnd.kinar' { Mime.application_vnd_kinar }
        'application/vnd.kde.kontour' { Mime.application_vnd_kde_kontour }
        'application/vnd.kde.kpresenter' { Mime.application_vnd_kde_kpresenter }
        'application/vnd.kde.kspread' { Mime.application_vnd_kde_kspread }
        'application/vnd.kahootz' { Mime.application_vnd_kahootz }
        'application/vnd.kde.kword' { Mime.application_vnd_kde_kword }
        'application/x-latex' { Mime.application_x_latex }
        'application/vnd.llamagraphics.life-balance.desktop' { Mime.application_vnd_llamagraphics_life_balance_desktop }
        'application/vnd.llamagraphics.life-balance.exchange+xml' { Mime.application_vnd_llamagraphics_life_balance_exchange_xml }
        'application/vnd.hhe.lesson-player' { Mime.application_vnd_hhe_lesson_player }
        'application/vnd.route66.link66+xml' { Mime.application_vnd_route66_link66_xml }
        'application/lost+xml' { Mime.application_lost_xml }
        'application/vnd.ms-lrm' { Mime.application_vnd_ms_lrm }
        'application/vnd.frogans.ltf' { Mime.application_vnd_frogans_ltf }
        'audio/vnd.lucent.voice' { Mime.audio_vnd_lucent_voice }
        'application/vnd.lotus-wordpro' { Mime.application_vnd_lotus_wordpro }
        'application/x-msmediaview' { Mime.application_x_msmediaview }
        'video/mpeg' { Mime.video_mpeg }
        'audio/mpeg' { Mime.audio_mpeg }
        'audio/x-mpegurl' { Mime.audio_x_mpegurl }
        'video/vnd.mpegurl' { Mime.video_vnd_mpegurl }
        'video/x-m4v' { Mime.video_x_m4v }
        'application/mathematica' { Mime.application_mathematica }
        'application/vnd.ecowin.chart' { Mime.application_vnd_ecowin_chart }
        'text/troff' { Mime.text_troff }
        'application/mathml+xml' { Mime.application_mathml_xml }
        'text/mathml' { Mime.text_mathml }
        'application/vnd.sqlite3' { Mime.application_vnd_sqlite3 }
        'application/vnd.mobius.mbk' { Mime.application_vnd_mobius_mbk }
        'application/mbox' { Mime.application_mbox }
        'application/vnd.medcalcdata' { Mime.application_vnd_medcalcdata }
        'application/vnd.mcd' { Mime.application_vnd_mcd }
        'text/vnd.curl.mcurl' { Mime.text_vnd_curl_mcurl }
        'application/x-msaccess' { Mime.application_x_msaccess }
        'image/vnd.ms-modi' { Mime.image_vnd_ms_modi }
        'model/mesh' { Mime.model_mesh }
        'application/vnd.mfmp' { Mime.application_vnd_mfmp }
        'application/vnd.proteus.magazine' { Mime.application_vnd_proteus_magazine }
        'application/vnd.mif' { Mime.application_vnd_mif }
        'video/mj2' { Mime.video_mj2 }
        'application/vnd.dolby.mlp' { Mime.application_vnd_dolby_mlp }
        'application/vnd.chipnuts.karaoke-mmd' { Mime.application_vnd_chipnuts_karaoke_mmd }
        'application/vnd.smaf' { Mime.application_vnd_smaf }
        'image/vnd.fujixerox.edmics-mmr' { Mime.image_vnd_fujixerox_edmics_mmr }
        'application/x-msmoney' { Mime.application_x_msmoney }
        'application/x-mobipocket-ebook' { Mime.application_x_mobipocket_ebook }
        'video/quicktime' { Mime.video_quicktime }
        'video/x-sgi-movie' { Mime.video_x_sgi_movie }
        'video/mp4' { Mime.video_mp4 }
        'application/x-iso9660-image' { Mime.application_x_iso9660_image }
        'application/yaml' { Mime.application_yaml }
        'application/mp4' { Mime.application_mp4 }
        'application/vnd.mophun.certificate' { Mime.application_vnd_mophun_certificate }
        'application/vnd.apple.installer+xml' { Mime.application_vnd_apple_installer_xml }
        'application/vnd.blueice.multipass' { Mime.application_vnd_blueice_multipass }
        'application/vnd.mophun.application' { Mime.application_vnd_mophun_application }
        'application/vnd.ms-project' { Mime.application_vnd_ms_project }
        'application/vnd.ibm.minipay' { Mime.application_vnd_ibm_minipay }
        'application/vnd.mobius.mqy' { Mime.application_vnd_mobius_mqy }
        'application/marc' { Mime.application_marc }
        'application/mediaservercontrol+xml' { Mime.application_mediaservercontrol_xml }
        'application/vnd.fdsn.mseed' { Mime.application_vnd_fdsn_mseed }
        'application/vnd.mseq' { Mime.application_vnd_mseq }
        'application/vnd.epson.msf' { Mime.application_vnd_epson_msf }
        'application/vnd.mobius.msl' { Mime.application_vnd_mobius_msl }
        'application/vnd.muvee.style' { Mime.application_vnd_muvee_style }
        'model/vnd.mts' { Mime.model_vnd_mts }
        'application/vnd.musician' { Mime.application_vnd_musician }
        'application/vnd.recordare.musicxml+xml' { Mime.application_vnd_recordare_musicxml_xml }
        'application/vnd.mfer' { Mime.application_vnd_mfer }
        'application/mxf' { Mime.application_mxf }
        'application/vnd.recordare.musicxml' { Mime.application_vnd_recordare_musicxml }
        'application/xv+xml' { Mime.application_xv_xml }
        'application/vnd.triscape.mxs' { Mime.application_vnd_triscape_mxs }
        'application/vnd.nokia.n-gage.symbian.install' { Mime.application_vnd_nokia_n_gage_symbian_install }
        'application/x-dtbncx+xml' { Mime.application_x_dtbncx_xml }
        'application/vnd.nokia.n-gage.data' { Mime.application_vnd_nokia_n_gage_data }
        'application/vnd.neurolanguage.nlu' { Mime.application_vnd_neurolanguage_nlu }
        'application/vnd.enliven' { Mime.application_vnd_enliven }
        'application/vnd.noblenet-directory' { Mime.application_vnd_noblenet_directory }
        'application/vnd.noblenet-sealer' { Mime.application_vnd_noblenet_sealer }
        'application/vnd.noblenet-web' { Mime.application_vnd_noblenet_web }
        'image/vnd.net-fpx' { Mime.image_vnd_net_fpx }
        'application/vnd.lotus-notes' { Mime.application_vnd_lotus_notes }
        'application/vnd.fujitsu.oasys2' { Mime.application_vnd_fujitsu_oasys2 }
        'application/vnd.fujitsu.oasys3' { Mime.application_vnd_fujitsu_oasys3 }
        'application/vnd.fujitsu.oasys' { Mime.application_vnd_fujitsu_oasys }
        'application/x-msbinder' { Mime.application_x_msbinder }
        'application/oda' { Mime.application_oda }
        'application/vnd.oasis.opendocument.database' { Mime.application_vnd_oasis_opendocument_database }
        'application/vnd.oasis.opendocument.chart' { Mime.application_vnd_oasis_opendocument_chart }
        'application/vnd.oasis.opendocument.formula' { Mime.application_vnd_oasis_opendocument_formula }
        'application/vnd.oasis.opendocument.formula-template' { Mime.application_vnd_oasis_opendocument_formula_template }
        'application/vnd.oasis.opendocument.graphics' { Mime.application_vnd_oasis_opendocument_graphics }
        'application/vnd.oasis.opendocument.image' { Mime.application_vnd_oasis_opendocument_image }
        'application/vnd.oasis.opendocument.presentation' { Mime.application_vnd_oasis_opendocument_presentation }
        'application/vnd.oasis.opendocument.spreadsheet' { Mime.application_vnd_oasis_opendocument_spreadsheet }
        'application/vnd.oasis.opendocument.text' { Mime.application_vnd_oasis_opendocument_text }
        'audio/ogg' { Mime.audio_ogg }
        'video/x-matroska' { Mime.video_x_matroska }
        'audio/x-matroska' { Mime.audio_x_matroska }
        'video/ogg' { Mime.video_ogg }
        'application/ogg' { Mime.application_ogg }
        'application/onenote' { Mime.application_onenote }
        'application/oebps-package+xml' { Mime.application_oebps_package_xml }
        'application/vnd.palm' { Mime.application_vnd_palm }
        'application/vnd.lotus-organizer' { Mime.application_vnd_lotus_organizer }
        'application/vnd.yamaha.openscoreformat' { Mime.application_vnd_yamaha_openscoreformat }
        'application/vnd.yamaha.openscoreformat.osfpvg+xml' { Mime.application_vnd_yamaha_openscoreformat_osfpvg_xml }
        'application/vnd.oasis.opendocument.chart-template' { Mime.application_vnd_oasis_opendocument_chart_template }
        'font/woff' { Mime.font_woff }
        'font/woff2' { Mime.font_woff2 }
        'application/x-redhat-package-manager' { Mime.application_x_redhat_package_manager }
        'application/x-perl' { Mime.application_x_perl }
        'audio/webm' { Mime.audio_webm }
        'video/webm' { Mime.video_webm }
        'image/webp' { Mime.image_webp }
        'application/x-font-otf' { Mime.application_x_font_otf }
        'font/otf' { Mime.font_otf }
        'application/vnd.oasis.opendocument.graphics-template' { Mime.application_vnd_oasis_opendocument_graphics_template }
        'application/vnd.oasis.opendocument.text-web' { Mime.application_vnd_oasis_opendocument_text_web }
        'application/vnd.oasis.opendocument.image-template' { Mime.application_vnd_oasis_opendocument_image_template }
        'application/vnd.oasis.opendocument.text-master' { Mime.application_vnd_oasis_opendocument_text_master }
        'application/vnd.oasis.opendocument.presentation-template' { Mime.application_vnd_oasis_opendocument_presentation_template }
        'application/vnd.oasis.opendocument.spreadsheet-template' { Mime.application_vnd_oasis_opendocument_spreadsheet_template }
        'application/vnd.oasis.opendocument.text-template' { Mime.application_vnd_oasis_opendocument_text_template }
        'application/vnd.openofficeorg.extension' { Mime.application_vnd_openofficeorg_extension }
        'text/x-pascal' { Mime.text_x_pascal }
        'application/pkcs10' { Mime.application_pkcs10 }
        'application/x-pkcs12' { Mime.application_x_pkcs12 }
        'application/x-pkcs7-certificates' { Mime.application_x_pkcs7_certificates }
        'application/pkcs7-mime' { Mime.application_pkcs7_mime }
        'application/x-pkcs7-certreqresp' { Mime.application_x_pkcs7_certreqresp }
        'application/pkcs7-signature' { Mime.application_pkcs7_signature }
        'application/vnd.powerbuilder6' { Mime.application_vnd_powerbuilder6 }
        'image/x-portable-bitmap' { Mime.image_x_portable_bitmap }
        'application/x-font-pcf' { Mime.application_x_font_pcf }
        'application/vnd.hp-pcl' { Mime.application_vnd_hp_pcl }
        'application/vnd.hp-pclxl' { Mime.application_vnd_hp_pclxl }
        'image/x-pict' { Mime.image_x_pict }
        'application/vnd.curl.pcurl' { Mime.application_vnd_curl_pcurl }
        'image/x-pcx' { Mime.image_x_pcx }
        'application/pdf' { Mime.application_pdf }
        'application/font-tdpfr' { Mime.application_font_tdpfr }
        'image/x-portable-graymap' { Mime.image_x_portable_graymap }
        'application/x-chess-pgn' { Mime.application_x_chess_pgn }
        'application/pgp-encrypted' { Mime.application_pgp_encrypted }
        'application/pkixcmp' { Mime.application_pkixcmp }
        'application/pkix-pkipath' { Mime.application_pkix_pkipath }
        'application/vnd.3gpp.pic-bw-large' { Mime.application_vnd_3gpp_pic_bw_large }
        'application/vnd.mobius.plc' { Mime.application_vnd_mobius_plc }
        'application/vnd.pocketlearn' { Mime.application_vnd_pocketlearn }
        'application/pls+xml' { Mime.application_pls_xml }
        'application/vnd.ctc-posml' { Mime.application_vnd_ctc_posml }
        'image/png' { Mime.image_png }
        'image/x-portable-anymap' { Mime.image_x_portable_anymap }
        'application/vnd.macports.portpkg' { Mime.application_vnd_macports_portpkg }
        'application/vnd.ms-powerpoint' { Mime.application_vnd_ms_powerpoint }
        'application/vnd.ms-powerpoint.template.macroenabled.12' { Mime.application_vnd_ms_powerpoint_template_macroenabled_12 }
        'application/vnd.openxmlformats-officedocument.presentationml.template' { Mime.application_vnd_openxmlformats_officedocument_presentationml_template }
        'application/vnd.ms-powerpoint.addin.macroenabled.12' { Mime.application_vnd_ms_powerpoint_addin_macroenabled_12 }
        'application/vnd.cups-ppd' { Mime.application_vnd_cups_ppd }
        'image/x-portable-pixmap' { Mime.image_x_portable_pixmap }
        'application/vnd.ms-powerpoint.slideshow.macroenabled.12' { Mime.application_vnd_ms_powerpoint_slideshow_macroenabled_12 }
        'application/vnd.openxmlformats-officedocument.presentationml.slideshow' { Mime.application_vnd_openxmlformats_officedocument_presentationml_slideshow }
        'application/vnd.ms-powerpoint.presentation.macroenabled.12' { Mime.application_vnd_ms_powerpoint_presentation_macroenabled_12 }
        'application/vnd.openxmlformats-officedocument.presentationml.presentation' { Mime.application_vnd_openxmlformats_officedocument_presentationml_presentation }
        'application/vnd.lotus-freelance' { Mime.application_vnd_lotus_freelance }
        'application/pics-rules' { Mime.application_pics_rules }
        'application/prql' { Mime.application_prql }
        'application/vnd.3gpp.pic-bw-small' { Mime.application_vnd_3gpp_pic_bw_small }
        'image/vnd.adobe.photoshop' { Mime.image_vnd_adobe_photoshop }
        'application/x-font-linux-psf' { Mime.application_x_font_linux_psf }
        'application/vnd.pvi.ptid1' { Mime.application_vnd_pvi_ptid1 }
        'application/x-mspublisher' { Mime.application_x_mspublisher }
        'application/vnd.3gpp.pic-bw-var' { Mime.application_vnd_3gpp_pic_bw_var }
        'application/vnd.3m.post-it-notes' { Mime.application_vnd_3m_post_it_notes }
        'text/x-python' { Mime.text_x_python }
        'audio/vnd.ms-playready.media.pya' { Mime.audio_vnd_ms_playready_media_pya }
        'video/vnd.ms-playready.media.pyv' { Mime.video_vnd_ms_playready_media_pyv }
        'application/vnd.epson.quickanime' { Mime.application_vnd_epson_quickanime }
        'application/vnd.intu.qbo' { Mime.application_vnd_intu_qbo }
        'application/vnd.intu.qfx' { Mime.application_vnd_intu_qfx }
        'application/vnd.publishare-delta-tree' { Mime.application_vnd_publishare_delta_tree }
        'application/vnd.quark.quarkxpress' { Mime.application_vnd_quark_quarkxpress }
        'audio/x-pn-realaudio' { Mime.audio_x_pn_realaudio }
        'application/vnd.rar' { Mime.application_vnd_rar }
        'application/x-rar-compressed' { Mime.application_x_rar_compressed }
        'image/x-cmu-raster' { Mime.image_x_cmu_raster }
        'application/vnd.ipunplugged.rcprofile' { Mime.application_vnd_ipunplugged_rcprofile }
        'application/rdf+xml' { Mime.application_rdf_xml }
        'application/vnd.data-vision.rdz' { Mime.application_vnd_data_vision_rdz }
        'application/vnd.businessobjects' { Mime.application_vnd_businessobjects }
        'application/x-dtbresource+xml' { Mime.application_x_dtbresource_xml }
        'image/x-rgb' { Mime.image_x_rgb }
        'application/reginfo+xml' { Mime.application_reginfo_xml }
        'application/resource-lists+xml' { Mime.application_resource_lists_xml }
        'image/vnd.fujixerox.edmics-rlc' { Mime.image_vnd_fujixerox_edmics_rlc }
        'application/resource-lists-diff+xml' { Mime.application_resource_lists_diff_xml }
        'application/vnd.rn-realmedia' { Mime.application_vnd_rn_realmedia }
        'audio/x-pn-realaudio-plugin' { Mime.audio_x_pn_realaudio_plugin }
        'application/vnd.jcp.javame.midlet-rms' { Mime.application_vnd_jcp_javame_midlet_rms }
        'application/relax-ng-compact-syntax' { Mime.application_relax_ng_compact_syntax }
        'application/x-rpm' { Mime.application_x_rpm }
        'application/vnd.nokia.radio-presets' { Mime.application_vnd_nokia_radio_presets }
        'application/vnd.nokia.radio-preset' { Mime.application_vnd_nokia_radio_preset }
        'application/sparql-query' { Mime.application_sparql_query }
        'application/rls-services+xml' { Mime.application_rls_services_xml }
        'application/rsd+xml' { Mime.application_rsd_xml }
        'application/rss+xml' { Mime.application_rss_xml }
        'application/rtf' { Mime.application_rtf }
        'text/richtext' { Mime.text_richtext }
        'application/vnd.yamaha.smaf-audio' { Mime.application_vnd_yamaha_smaf_audio }
        'application/sbml+xml' { Mime.application_sbml_xml }
        'application/vnd.ibm.secure-container' { Mime.application_vnd_ibm_secure_container }
        'application/x-msschedule' { Mime.application_x_msschedule }
        'application/vnd.lotus-screencam' { Mime.application_vnd_lotus_screencam }
        'application/scvp-cv-request' { Mime.application_scvp_cv_request }
        'application/scvp-cv-response' { Mime.application_scvp_cv_response }
        'text/vnd.curl.scurl' { Mime.text_vnd_curl_scurl }
        'application/vnd.stardivision.draw' { Mime.application_vnd_stardivision_draw }
        'application/vnd.stardivision.calc' { Mime.application_vnd_stardivision_calc }
        'application/vnd.stardivision.impress' { Mime.application_vnd_stardivision_impress }
        'application/vnd.solent.sdkm+xml' { Mime.application_vnd_solent_sdkm_xml }
        'application/sdp' { Mime.application_sdp }
        'application/vnd.stardivision.writer' { Mime.application_vnd_stardivision_writer }
        'application/vnd.seemail' { Mime.application_vnd_seemail }
        'application/vnd.sema' { Mime.application_vnd_sema }
        'application/vnd.semd' { Mime.application_vnd_semd }
        'application/vnd.semf' { Mime.application_vnd_semf }
        'application/java-serialized-object' { Mime.application_java_serialized_object }
        'application/set-payment-initiation' { Mime.application_set_payment_initiation }
        'application/set-registration-initiation' { Mime.application_set_registration_initiation }
        'application/vnd.hydrostatix.sof-data' { Mime.application_vnd_hydrostatix_sof_data }
        'application/vnd.spotfire.sfs' { Mime.application_vnd_spotfire_sfs }
        'application/vnd.stardivision.writer-global' { Mime.application_vnd_stardivision_writer_global }
        'text/sgml' { Mime.text_sgml }
        'application/x-sh' { Mime.application_x_sh }
        'application/x-shar' { Mime.application_x_shar }
        'application/shf+xml' { Mime.application_shf_xml }
        'text/vnd.wap.si' { Mime.text_vnd_wap_si }
        'application/vnd.wap.sic' { Mime.application_vnd_wap_sic }
        'application/vnd.symbian.install' { Mime.application_vnd_symbian_install }
        'application/x-stuffit' { Mime.application_x_stuffit }
        'application/x-stuffitx' { Mime.application_x_stuffitx }
        'application/vnd.koan' { Mime.application_vnd_koan }
        'text/vnd.wap.sl' { Mime.text_vnd_wap_sl }
        'application/vnd.wap.slc' { Mime.application_vnd_wap_slc }
        'application/vnd.ms-powerpoint.slide.macroenabled.12' { Mime.application_vnd_ms_powerpoint_slide_macroenabled_12 }
        'application/vnd.openxmlformats-officedocument.presentationml.slide' { Mime.application_vnd_openxmlformats_officedocument_presentationml_slide }
        'application/vnd.epson.salt' { Mime.application_vnd_epson_salt }
        'application/vnd.stardivision.math' { Mime.application_vnd_stardivision_math }
        'application/smil+xml' { Mime.application_smil_xml }
        'application/x-font-snf' { Mime.application_x_font_snf }
        'application/vnd.yamaha.smaf-phrase' { Mime.application_vnd_yamaha_smaf_phrase }
        'application/x-futuresplash' { Mime.application_x_futuresplash }
        'text/vnd.in3d.spot' { Mime.text_vnd_in3d_spot }
        'application/scvp-vp-response' { Mime.application_scvp_vp_response }
        'application/scvp-vp-request' { Mime.application_scvp_vp_request }
        'application/x-wais-source' { Mime.application_x_wais_source }
        'application/sparql-results+xml' { Mime.application_sparql_results_xml }
        'application/vnd.kodak-descriptor' { Mime.application_vnd_kodak_descriptor }
        'application/vnd.epson.ssf' { Mime.application_vnd_epson_ssf }
        'application/ssml+xml' { Mime.application_ssml_xml }
        'application/vnd.sun.xml.calc.template' { Mime.application_vnd_sun_xml_calc_template }
        'application/vnd.sun.xml.draw.template' { Mime.application_vnd_sun_xml_draw_template }
        'application/vnd.wt.stf' { Mime.application_vnd_wt_stf }
        'application/vnd.sun.xml.impress.template' { Mime.application_vnd_sun_xml_impress_template }
        'application/hyperstudio' { Mime.application_hyperstudio }
        'application/vnd.ms-pki.stl' { Mime.application_vnd_ms_pki_stl }
        'application/vnd.pg.format' { Mime.application_vnd_pg_format }
        'application/vnd.sun.xml.writer.template' { Mime.application_vnd_sun_xml_writer_template }
        'application/vnd.sus-calendar' { Mime.application_vnd_sus_calendar }
        'application/x-sv4cpio' { Mime.application_x_sv4cpio }
        'application/x-sv4crc' { Mime.application_x_sv4crc }
        'application/vnd.svd' { Mime.application_vnd_svd }
        'image/svg+xml' { Mime.image_svg_xml }
        'application/x-shockwave-flash' { Mime.application_x_shockwave_flash }
        'application/vnd.arastra.swi' { Mime.application_vnd_arastra_swi }
        'application/vnd.sun.xml.calc' { Mime.application_vnd_sun_xml_calc }
        'application/vnd.sun.xml.draw' { Mime.application_vnd_sun_xml_draw }
        'application/vnd.sun.xml.writer.global' { Mime.application_vnd_sun_xml_writer_global }
        'application/vnd.sun.xml.impress' { Mime.application_vnd_sun_xml_impress }
        'application/vnd.sun.xml.math' { Mime.application_vnd_sun_xml_math }
        'application/vnd.sun.xml.writer' { Mime.application_vnd_sun_xml_writer }
        'application/vnd.tao.intent-module-archive' { Mime.application_vnd_tao_intent_module_archive }
        'application/x-tar' { Mime.application_x_tar }
        'application/vnd.3gpp2.tcap' { Mime.application_vnd_3gpp2_tcap }
        'application/x-tcl' { Mime.application_x_tcl }
        'application/vnd.smart.teacher' { Mime.application_vnd_smart_teacher }
        'application/x-tex' { Mime.application_x_tex }
        'application/x-texinfo' { Mime.application_x_texinfo }
        'application/x-tex-tfm' { Mime.application_x_tex_tfm }
        'image/tiff' { Mime.image_tiff }
        'application/vnd.tmobile-livetv' { Mime.application_vnd_tmobile_livetv }
        'application/x-bittorrent' { Mime.application_x_bittorrent }
        'application/vnd.groove-tool-template' { Mime.application_vnd_groove_tool_template }
        'application/vnd.trid.tpt' { Mime.application_vnd_trid_tpt }
        'application/vnd.trueapp' { Mime.application_vnd_trueapp }
        'application/x-msterminal' { Mime.application_x_msterminal }
        'text/tab-separated-values' { Mime.text_tab_separated_values }
        'application/x-font-ttf' { Mime.application_x_font_ttf }
        'application/vnd.simtech-mindmapper' { Mime.application_vnd_simtech_mindmapper }
        'application/vnd.genomatix.tuxedo' { Mime.application_vnd_genomatix_tuxedo }
        'application/vnd.mobius.txf' { Mime.application_vnd_mobius_txf }
        'application/vnd.ufdl' { Mime.application_vnd_ufdl }
        'test/mimetype' { Mime.test_mimetype }
        'application/vnd.umajin' { Mime.application_vnd_umajin }
        'application/vnd.unity' { Mime.application_vnd_unity }
        'application/vnd.uoml+xml' { Mime.application_vnd_uoml_xml }
        'text/uri-list' { Mime.text_uri_list }
        'application/x-ustar' { Mime.application_x_ustar }
        'application/vnd.uiq.theme' { Mime.application_vnd_uiq_theme }
        'text/x-uuencode' { Mime.text_x_uuencode }
        'application/x-cdlink' { Mime.application_x_cdlink }
        'text/x-vcard' { Mime.text_x_vcard }
        'application/vnd.groove-vcard' { Mime.application_vnd_groove_vcard }
        'text/x-vcalendar' { Mime.text_x_vcalendar }
        'application/vnd.vcx' { Mime.application_vnd_vcx }
        'application/vnd.visionary' { Mime.application_vnd_visionary }
        'video/vnd.vivo' { Mime.video_vnd_vivo }
        'model/vrml' { Mime.model_vrml }
        'application/vnd.visio' { Mime.application_vnd_visio }
        'application/vnd.vsf' { Mime.application_vnd_vsf }
        'model/vnd.vtu' { Mime.model_vnd_vtu }
        'application/voicexml+xml' { Mime.application_voicexml_xml }
        'application/x-doom' { Mime.application_x_doom }
        'video/mp2t' { Mime.video_mp2t }
        'audio/vnd.wav' { Mime.audio_vnd_wav }
        'audio/x-ms-wax' { Mime.audio_x_ms_wax }
        'image/vnd.wap.wbmp' { Mime.image_vnd_wap_wbmp }
        'application/vnd.criticaltools.wbs+xml' { Mime.application_vnd_criticaltools_wbs_xml }
        'application/vnd.wap.wbxml' { Mime.application_vnd_wap_wbxml }
        'application/vnd.ms-works' { Mime.application_vnd_ms_works }
        'video/x-ms-wm' { Mime.video_x_ms_wm }
        'audio/x-ms-wma' { Mime.audio_x_ms_wma }
        'application/x-ms-wmd' { Mime.application_x_ms_wmd }
        'application/x-msmetafile' { Mime.application_x_msmetafile }
        'text/vnd.wap.wml' { Mime.text_vnd_wap_wml }
        'application/vnd.wap.wmlc' { Mime.application_vnd_wap_wmlc }
        'text/vnd.wap.wmlscript' { Mime.text_vnd_wap_wmlscript }
        'application/vnd.wap.wmlscriptc' { Mime.application_vnd_wap_wmlscriptc }
        'video/x-ms-wmv' { Mime.video_x_ms_wmv }
        'video/x-ms-wmx' { Mime.video_x_ms_wmx }
        'application/x-ms-wmz' { Mime.application_x_ms_wmz }
        'application/vnd.wordperfect' { Mime.application_vnd_wordperfect }
        'application/vnd.ms-wpl' { Mime.application_vnd_ms_wpl }
        'application/vnd.wqd' { Mime.application_vnd_wqd }
        'application/x-mswrite' { Mime.application_x_mswrite }
        'application/wsdl+xml' { Mime.application_wsdl_xml }
        'application/wspolicy+xml' { Mime.application_wspolicy_xml }
        'application/vnd.webturbo' { Mime.application_vnd_webturbo }
        'video/x-ms-wvx' { Mime.video_x_ms_wvx }
        'application/vnd.hzn-3d-crossword' { Mime.application_vnd_hzn_3d_crossword }
        'application/x-silverlight-app' { Mime.application_x_silverlight_app }
        'application/vnd.xara' { Mime.application_vnd_xara }
        'application/x-ms-xbap' { Mime.application_x_ms_xbap }
        'application/vnd.fujixerox.docuworks.binder' { Mime.application_vnd_fujixerox_docuworks_binder }
        'image/x-xbitmap' { Mime.image_x_xbitmap }
        'application/vnd.syncml.dm+xml' { Mime.application_vnd_syncml_dm_xml }
        'application/vnd.adobe.xdp+xml' { Mime.application_vnd_adobe_xdp_xml }
        'application/vnd.fujixerox.docuworks' { Mime.application_vnd_fujixerox_docuworks }
        'application/xenc+xml' { Mime.application_xenc_xml }
        'application/patch-ops-error+xml' { Mime.application_patch_ops_error_xml }
        'application/vnd.adobe.xfdf' { Mime.application_vnd_adobe_xfdf }
        'application/vnd.xfdl' { Mime.application_vnd_xfdl }
        'application/xhtml+xml' { Mime.application_xhtml_xml }
        'image/vnd.xiff' { Mime.image_vnd_xiff }
        'application/vnd.ms-excel' { Mime.application_vnd_ms_excel }
        'application/vnd.ms-excel.addin.macroenabled.12' { Mime.application_vnd_ms_excel_addin_macroenabled_12 }
        'application/vnd.ms-excel.sheet.binary.macroenabled.12' { Mime.application_vnd_ms_excel_sheet_binary_macroenabled_12 }
        'application/vnd.ms-excel.sheet.macroenabled.12' { Mime.application_vnd_ms_excel_sheet_macroenabled_12 }
        'application/vnd.openxmlformats-officedocument.spreadsheetml.sheet' { Mime.application_vnd_openxmlformats_officedocument_spreadsheetml_sheet }
        'application/vnd.ms-excel.template.macroenabled.12' { Mime.application_vnd_ms_excel_template_macroenabled_12 }
        'application/vnd.openxmlformats-officedocument.spreadsheetml.template' { Mime.application_vnd_openxmlformats_officedocument_spreadsheetml_template }
        'application/xml' { Mime.application_xml }
        'application/vnd.olpc-sugar' { Mime.application_vnd_olpc_sugar }
        'application/xop+xml' { Mime.application_xop_xml }
        'application/x-xpinstall' { Mime.application_x_xpinstall }
        'image/x-xpixmap' { Mime.image_x_xpixmap }
        'application/vnd.is-xpr' { Mime.application_vnd_is_xpr }
        'application/vnd.ms-xpsdocument' { Mime.application_vnd_ms_xpsdocument }
        'application/vnd.intercon.formnet' { Mime.application_vnd_intercon_formnet }
        'application/xslt+xml' { Mime.application_xslt_xml }
        'application/vnd.syncml+xml' { Mime.application_vnd_syncml_xml }
        'application/xspf+xml' { Mime.application_xspf_xml }
        'application/vnd.mozilla.xul+xml' { Mime.application_vnd_mozilla_xul_xml }
        'image/x-xwindowdump' { Mime.image_x_xwindowdump }
        'chemical/x-xyz' { Mime.chemical_x_xyz }
        'application/vnd.zzazz.deck+xml' { Mime.application_vnd_zzazz_deck_xml }
        'application/zip' { Mime.application_zip }
        'application/x-zip-compressed' { Mime.application_x_zip_compressed }
        'application/zip-compressed' { Mime.application_zip_compressed }
        'application/vnd.zul' { Mime.application_vnd_zul }
        'application/vnd.handheld-entertainment+xml' { Mime.application_vnd_handheld_entertainment_xml }
        'image/x-adobe-dng' { Mime.image_x_adobe_dng }
        'image/x-sony-arw' { Mime.image_x_sony_arw }
        'image/x-canon-cr2' { Mime.image_x_canon_cr2 }
        'image/x-canon-crw' { Mime.image_x_canon_crw }
        'image/x-kodak-dcr' { Mime.image_x_kodak_dcr }
        'image/x-epson-erf' { Mime.image_x_epson_erf }
        'image/x-kodak-k25' { Mime.image_x_kodak_k25 }
        'image/x-kodak-kdc' { Mime.image_x_kodak_kdc }
        'image/x-minolta-mrw' { Mime.image_x_minolta_mrw }
        'image/x-nikon-nef' { Mime.image_x_nikon_nef }
        'image/x-olympus-orf' { Mime.image_x_olympus_orf }
        'image/x-pentax-pef' { Mime.image_x_pentax_pef }
        'image/x-fuji-raf' { Mime.image_x_fuji_raf }
        'image/x-panasonic-raw' { Mime.image_x_panasonic_raw }
        'audio/flac' { Mime.audio_flac }
        'image/x-sony-sr2' { Mime.image_x_sony_sr2 }
        'image/x-sony-srf' { Mime.image_x_sony_srf }
        'image/x-sigma-x3f' { Mime.image_x_sigma_x3f }
        else { none }
    }
}
