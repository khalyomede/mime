module mime

pub enum Mime {
    text_html
    application_json
}
