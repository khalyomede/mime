module mime

pub fn (m Mime) str() string {
    return match m {
        .application_vnd_lotus_1_2_3 { 'application/vnd.lotus-1-2-3' }
        .text_vnd_in3d_3dml { 'text/vnd.in3d.3dml' }
        .video_3gpp2 { 'video/3gpp2' }
        .image_avif { 'image/avif' }
        .image_avif_sequence { 'image/avif-sequence' }
        .application_x_krita { 'application/x-krita' }
        .image_heic { 'image/heic' }
        .video_3gpp { 'video/3gpp' }
        .audio_3gpp2 { 'audio/3gpp2' }
        .application_x_7z_compressed { 'application/x-7z-compressed' }
        .application_octet_stream { 'application/octet-stream' }
        .application_x_authorware_bin { 'application/x-authorware-bin' }
        .image_x_icns { 'image/x-icns' }
        .audio_mp4 { 'audio/mp4' }
        .audio_aac { 'audio/aac' }
        .audio_mp4a_latm { 'audio/mp4a-latm' }
        .audio_aacp { 'audio/aacp' }
        .application_x_authorware_map { 'application/x-authorware-map' }
        .application_x_authorware_seg { 'application/x-authorware-seg' }
        .application_x_abiword { 'application/x-abiword' }
        .application_vnd_americandynamics_acc { 'application/vnd.americandynamics.acc' }
        .application_x_ace_compressed { 'application/x-ace-compressed' }
        .application_vnd_acucobol { 'application/vnd.acucobol' }
        .application_vnd_acucorp { 'application/vnd.acucorp' }
        .audio_adpcm { 'audio/adpcm' }
        .application_vnd_audiograph { 'application/vnd.audiograph' }
        .application_x_font_type1 { 'application/x-font-type1' }
        .application_vnd_ibm_modcap { 'application/vnd.ibm.modcap' }
        .application_postscript { 'application/postscript' }
        .application_vnd_adobe_air_application_installer_package_zip { 'application/vnd.adobe.air-application-installer-package+zip' }
        .application_vnd_amiga_ami { 'application/vnd.amiga.ami' }
        .application_vnd_android_package_archive { 'application/vnd.android.package-archive' }
        .application_x_ms_application { 'application/x-ms-application' }
        .application_vnd_lotus_approach { 'application/vnd.lotus-approach' }
        .application_pgp_signature { 'application/pgp-signature' }
        .video_x_ms_asf { 'video/x-ms-asf' }
        .text_x_asm { 'text/x-asm' }
        .application_vnd_accpac_simply_aso { 'application/vnd.accpac.simply.aso' }
        .application_atom_xml { 'application/atom+xml' }
        .application_atomcat_xml { 'application/atomcat+xml' }
        .application_atomsvc_xml { 'application/atomsvc+xml' }
        .application_vnd_antix_game_component { 'application/vnd.antix.game-component' }
        .audio_basic { 'audio/basic' }
        .video_x_msvideo { 'video/x-msvideo' }
        .application_applixware { 'application/applixware' }
        .application_vnd_airzip_filesecure_azf { 'application/vnd.airzip.filesecure.azf' }
        .application_vnd_airzip_filesecure_azs { 'application/vnd.airzip.filesecure.azs' }
        .application_vnd_amazon_ebook { 'application/vnd.amazon.ebook' }
        .application_x_msdownload { 'application/x-msdownload' }
        .application_x_bcpio { 'application/x-bcpio' }
        .application_x_font_bdf { 'application/x-font-bdf' }
        .application_vnd_syncml_dm_wbxml { 'application/vnd.syncml.dm+wbxml' }
        .application_vnd_fujitsu_oasysprs { 'application/vnd.fujitsu.oasysprs' }
        .application_vnd_bmi { 'application/vnd.bmi' }
        .image_bmp { 'image/bmp' }
        .application_vnd_framemaker { 'application/vnd.framemaker' }
        .application_vnd_previewsystems_box { 'application/vnd.previewsystems.box' }
        .application_x_bzip2 { 'application/x-bzip2' }
        .image_prs_btif { 'image/prs.btif' }
        .application_x_bzip { 'application/x-bzip' }
        .text_x_c { 'text/x-c' }
        .application_vnd_clonk_c4group { 'application/vnd.clonk.c4group' }
        .application_vnd_ms_cab_compressed { 'application/vnd.ms-cab-compressed' }
        .application_vnd_curl_car { 'application/vnd.curl.car' }
        .application_vnd_ms_pki_seccat { 'application/vnd.ms-pki.seccat' }
        .application_x_director { 'application/x-director' }
        .application_ccxml_xml { 'application/ccxml+xml' }
        .application_vnd_contact_cmsg { 'application/vnd.contact.cmsg' }
        .application_x_netcdf { 'application/x-netcdf' }
        .application_vnd_mediastation_cdkey { 'application/vnd.mediastation.cdkey' }
        .chemical_x_cdx { 'chemical/x-cdx' }
        .application_vnd_chemdraw_xml { 'application/vnd.chemdraw+xml' }
        .application_vnd_cinderella { 'application/vnd.cinderella' }
        .application_pkix_cert { 'application/pkix-cert' }
        .image_cgm { 'image/cgm' }
        .application_x_chat { 'application/x-chat' }
        .application_vnd_ms_htmlhelp { 'application/vnd.ms-htmlhelp' }
        .application_vnd_kde_kchart { 'application/vnd.kde.kchart' }
        .chemical_x_cif { 'chemical/x-cif' }
        .application_vnd_anser_web_certificate_issue_initiation { 'application/vnd.anser-web-certificate-issue-initiation' }
        .application_vnd_ms_artgalry { 'application/vnd.ms-artgalry' }
        .application_vnd_claymore { 'application/vnd.claymore' }
        .application_java_vm { 'application/java-vm' }
        .application_vnd_crick_clicker_keyboard { 'application/vnd.crick.clicker.keyboard' }
        .application_vnd_crick_clicker_palette { 'application/vnd.crick.clicker.palette' }
        .application_vnd_crick_clicker_template { 'application/vnd.crick.clicker.template' }
        .application_vnd_crick_clicker_wordbank { 'application/vnd.crick.clicker.wordbank' }
        .application_vnd_crick_clicker { 'application/vnd.crick.clicker' }
        .application_x_msclip { 'application/x-msclip' }
        .application_vnd_cosmocaller { 'application/vnd.cosmocaller' }
        .chemical_x_cmdf { 'chemical/x-cmdf' }
        .chemical_x_cml { 'chemical/x-cml' }
        .application_vnd_yellowriver_custom_menu { 'application/vnd.yellowriver-custom-menu' }
        .image_x_cmx { 'image/x-cmx' }
        .application_vnd_rim_cod { 'application/vnd.rim.cod' }
        .text_plain { 'text/plain' }
        .application_vnd_debian_binary_package { 'application/vnd.debian.binary-package' }
        .text_markdown { 'text/markdown' }
        .application_wasm { 'application/wasm' }
        .application_x_cpio { 'application/x-cpio' }
        .application_mac_compactpro { 'application/mac-compactpro' }
        .application_x_mscardfile { 'application/x-mscardfile' }
        .application_pkix_crl { 'application/pkix-crl' }
        .application_x_x509_ca_cert { 'application/x-x509-ca-cert' }
        .application_x_csh { 'application/x-csh' }
        .chemical_x_csml { 'chemical/x-csml' }
        .application_vnd_commonspace { 'application/vnd.commonspace' }
        .text_css { 'text/css' }
        .text_csv { 'text/csv' }
        .application_cu_seeme { 'application/cu-seeme' }
        .text_vnd_curl { 'text/vnd.curl' }
        .application_prs_cww { 'application/prs.cww' }
        .application_vnd_mobius_daf { 'application/vnd.mobius.daf' }
        .application_vnd_fdsn_seed { 'application/vnd.fdsn.seed' }
        .application_davmount_xml { 'application/davmount+xml' }
        .text_vnd_curl_dcurl { 'text/vnd.curl.dcurl' }
        .application_vnd_oma_dd2_xml { 'application/vnd.oma.dd2+xml' }
        .application_vnd_fujixerox_ddd { 'application/vnd.fujixerox.ddd' }
        .application_x_debian_package { 'application/x-debian-package' }
        .application_vnd_dreamfactory { 'application/vnd.dreamfactory' }
        .application_vnd_mobius_dis { 'application/vnd.mobius.dis' }
        .image_vnd_djvu { 'image/vnd.djvu' }
        .application_vnd_dna { 'application/vnd.dna' }
        .application_msword { 'application/msword' }
        .application_vnd_ms_word_document_macroenabled_12 { 'application/vnd.ms-word.document.macroenabled.12' }
        .application_vnd_openxmlformats_officedocument_wordprocessingml_document { 'application/vnd.openxmlformats-officedocument.wordprocessingml.document' }
        .application_vnd_ms_word_template_macroenabled_12 { 'application/vnd.ms-word.template.macroenabled.12' }
        .application_vnd_openxmlformats_officedocument_wordprocessingml_template { 'application/vnd.openxmlformats-officedocument.wordprocessingml.template' }
        .application_vnd_osgi_dp { 'application/vnd.osgi.dp' }
        .application_vnd_dpgraph { 'application/vnd.dpgraph' }
        .text_prs_lines_tag { 'text/prs.lines.tag' }
        .application_x_dtbook_xml { 'application/x-dtbook+xml' }
        .application_xml_dtd { 'application/xml-dtd' }
        .audio_vnd_dts { 'audio/vnd.dts' }
        .audio_vnd_dts_hd { 'audio/vnd.dts.hd' }
        .application_x_dvi { 'application/x-dvi' }
        .model_vnd_dwf { 'model/vnd.dwf' }
        .image_vnd_dwg { 'image/vnd.dwg' }
        .image_vnd_dxf { 'image/vnd.dxf' }
        .application_vnd_spotfire_dxp { 'application/vnd.spotfire.dxp' }
        .audio_vnd_nuera_ecelp4800 { 'audio/vnd.nuera.ecelp4800' }
        .audio_vnd_nuera_ecelp7470 { 'audio/vnd.nuera.ecelp7470' }
        .audio_vnd_nuera_ecelp9600 { 'audio/vnd.nuera.ecelp9600' }
        .application_ecmascript { 'application/ecmascript' }
        .application_vnd_novadigm_edm { 'application/vnd.novadigm.edm' }
        .application_vnd_novadigm_edx { 'application/vnd.novadigm.edx' }
        .application_vnd_picsel { 'application/vnd.picsel' }
        .application_vnd_pg_osasli { 'application/vnd.pg.osasli' }
        .message_rfc822 { 'message/rfc822' }
        .application_emma_xml { 'application/emma+xml' }
        .audio_vnd_digital_winds { 'audio/vnd.digital-winds' }
        .application_vnd_ms_fontobject { 'application/vnd.ms-fontobject' }
        .application_epub_zip { 'application/epub+zip' }
        .application_vnd_eszigno3_xml { 'application/vnd.eszigno3+xml' }
        .application_vnd_epson_esf { 'application/vnd.epson.esf' }
        .text_x_setext { 'text/x-setext' }
        .application_vnd_novadigm_ext { 'application/vnd.novadigm.ext' }
        .application_andrew_inset { 'application/andrew-inset' }
        .application_vnd_ezpix_album { 'application/vnd.ezpix-album' }
        .application_vnd_ezpix_package { 'application/vnd.ezpix-package' }
        .text_x_fortran { 'text/x-fortran' }
        .video_x_f4v { 'video/x-f4v' }
        .image_vnd_fastbidsheet { 'image/vnd.fastbidsheet' }
        .application_vnd_fdf { 'application/vnd.fdf' }
        .application_vnd_denovo_fcselayout_link { 'application/vnd.denovo.fcselayout-link' }
        .application_vnd_fujitsu_oasysgp { 'application/vnd.fujitsu.oasysgp' }
        .image_x_freehand { 'image/x-freehand' }
        .application_x_xfig { 'application/x-xfig' }
        .video_x_fli { 'video/x-fli' }
        .application_vnd_micrografx_flo { 'application/vnd.micrografx.flo' }
        .video_x_flv { 'video/x-flv' }
        .application_vnd_kde_kivio { 'application/vnd.kde.kivio' }
        .text_vnd_fmi_flexstor { 'text/vnd.fmi.flexstor' }
        .text_vnd_fly { 'text/vnd.fly' }
        .application_vnd_frogans_fnc { 'application/vnd.frogans.fnc' }
        .image_vnd_fpx { 'image/vnd.fpx' }
        .application_vnd_fsc_weblaunch { 'application/vnd.fsc.weblaunch' }
        .image_vnd_fst { 'image/vnd.fst' }
        .application_vnd_fluxtime_clip { 'application/vnd.fluxtime.clip' }
        .application_vnd_anser_web_funds_transfer_initiation { 'application/vnd.anser-web-funds-transfer-initiation' }
        .video_vnd_fvt { 'video/vnd.fvt' }
        .application_vnd_fuzzysheet { 'application/vnd.fuzzysheet' }
        .image_g3fax { 'image/g3fax' }
        .application_vnd_groove_account { 'application/vnd.groove-account' }
        .model_vnd_gdl { 'model/vnd.gdl' }
        .application_vnd_dynageo { 'application/vnd.dynageo' }
        .application_vnd_geometry_explorer { 'application/vnd.geometry-explorer' }
        .application_vnd_geogebra_file { 'application/vnd.geogebra.file' }
        .application_vnd_geogebra_tool { 'application/vnd.geogebra.tool' }
        .application_vnd_groove_help { 'application/vnd.groove-help' }
        .image_gif { 'image/gif' }
        .application_vnd_groove_identity_message { 'application/vnd.groove-identity-message' }
        .application_vnd_gmx { 'application/vnd.gmx' }
        .application_x_gnumeric { 'application/x-gnumeric' }
        .application_vnd_flographit { 'application/vnd.flographit' }
        .application_vnd_grafeq { 'application/vnd.grafeq' }
        .application_srgs { 'application/srgs' }
        .application_vnd_groove_injector { 'application/vnd.groove-injector' }
        .application_srgs_xml { 'application/srgs+xml' }
        .application_x_font_ghostscript { 'application/x-font-ghostscript' }
        .application_x_gtar { 'application/x-gtar' }
        .application_vnd_groove_tool_message { 'application/vnd.groove-tool-message' }
        .model_vnd_gtw { 'model/vnd.gtw' }
        .text_vnd_graphviz { 'text/vnd.graphviz' }
        .application_x_gzip { 'application/x-gzip' }
        .application_gzip { 'application/gzip' }
        .video_h261 { 'video/h261' }
        .gcode { 'gcode' }
        .video_h263 { 'video/h263' }
        .video_h264 { 'video/h264' }
        .application_vnd_hbci { 'application/vnd.hbci' }
        .application_vnd_gerber { 'application/vnd.gerber' }
        .application_x_hdf { 'application/x-hdf' }
        .application_winhlp { 'application/winhlp' }
        .application_vnd_hp_hpgl { 'application/vnd.hp-hpgl' }
        .application_vnd_hp_hpid { 'application/vnd.hp-hpid' }
        .application_vnd_hp_hps { 'application/vnd.hp-hps' }
        .application_mac_binhex40 { 'application/mac-binhex40' }
        .application_vnd_kenameaapp { 'application/vnd.kenameaapp' }
        .text_html { 'text/html' }
        .application_vnd_yamaha_hv_dic { 'application/vnd.yamaha.hv-dic' }
        .application_vnd_yamaha_hv_voice { 'application/vnd.yamaha.hv-voice' }
        .application_vnd_yamaha_hv_script { 'application/vnd.yamaha.hv-script' }
        .application_vnd_iccprofile { 'application/vnd.iccprofile' }
        .x_conference_x_cooltalk { 'x-conference/x-cooltalk' }
        .image_x_icon { 'image/x-icon' }
        .text_calendar { 'text/calendar' }
        .image_ief { 'image/ief' }
        .application_vnd_shana_informed_formdata { 'application/vnd.shana.informed.formdata' }
        .model_iges { 'model/iges' }
        .application_vnd_igloader { 'application/vnd.igloader' }
        .application_vnd_micrografx_igx { 'application/vnd.micrografx.igx' }
        .application_vnd_shana_informed_interchange { 'application/vnd.shana.informed.interchange' }
        .application_vnd_accpac_simply_imp { 'application/vnd.accpac.simply.imp' }
        .application_vnd_ms_ims { 'application/vnd.ms-ims' }
        .application_vnd_shana_informed_package { 'application/vnd.shana.informed.package' }
        .application_vnd_ibm_rights_management { 'application/vnd.ibm.rights-management' }
        .application_vnd_irepository_package_xml { 'application/vnd.irepository.package+xml' }
        .application_vnd_shana_informed_formtemplate { 'application/vnd.shana.informed.formtemplate' }
        .application_vnd_immervision_ivp { 'application/vnd.immervision-ivp' }
        .application_vnd_immervision_ivu { 'application/vnd.immervision-ivu' }
        .text_vnd_sun_j2me_app_descriptor { 'text/vnd.sun.j2me.app-descriptor' }
        .application_vnd_jam { 'application/vnd.jam' }
        .application_java_archive { 'application/java-archive' }
        .text_x_java_source { 'text/x-java-source' }
        .application_vnd_jisp { 'application/vnd.jisp' }
        .application_vnd_hp_jlyt { 'application/vnd.hp-jlyt' }
        .application_x_java_jnlp_file { 'application/x-java-jnlp-file' }
        .application_vnd_joost_joda_archive { 'application/vnd.joost.joda-archive' }
        .image_jpeg { 'image/jpeg' }
        .image_pjpeg { 'image/pjpeg' }
        .video_jpm { 'video/jpm' }
        .video_jpeg { 'video/jpeg' }
        .application_x_trash { 'application/x-trash' }
        .application_x_shellscript { 'application/x-shellscript' }
        .text_javascript { 'text/javascript' }
        .application_json { 'application/json' }
        .audio_midi { 'audio/midi' }
        .audio_aiff { 'audio/aiff' }
        .audio_opus { 'audio/opus' }
        .application_vnd_kde_karbon { 'application/vnd.kde.karbon' }
        .application_vnd_kde_kformula { 'application/vnd.kde.kformula' }
        .application_vnd_kidspiration { 'application/vnd.kidspiration' }
        .application_x_killustrator { 'application/x-killustrator' }
        .application_vnd_google_earth_kml_xml { 'application/vnd.google-earth.kml+xml' }
        .application_vnd_google_earth_kmz { 'application/vnd.google-earth.kmz' }
        .application_vnd_kinar { 'application/vnd.kinar' }
        .application_vnd_kde_kontour { 'application/vnd.kde.kontour' }
        .application_vnd_kde_kpresenter { 'application/vnd.kde.kpresenter' }
        .application_vnd_kde_kspread { 'application/vnd.kde.kspread' }
        .application_vnd_kahootz { 'application/vnd.kahootz' }
        .application_vnd_kde_kword { 'application/vnd.kde.kword' }
        .application_x_latex { 'application/x-latex' }
        .application_vnd_llamagraphics_life_balance_desktop { 'application/vnd.llamagraphics.life-balance.desktop' }
        .application_vnd_llamagraphics_life_balance_exchange_xml { 'application/vnd.llamagraphics.life-balance.exchange+xml' }
        .application_vnd_hhe_lesson_player { 'application/vnd.hhe.lesson-player' }
        .application_vnd_route66_link66_xml { 'application/vnd.route66.link66+xml' }
        .application_lost_xml { 'application/lost+xml' }
        .application_vnd_ms_lrm { 'application/vnd.ms-lrm' }
        .application_vnd_frogans_ltf { 'application/vnd.frogans.ltf' }
        .audio_vnd_lucent_voice { 'audio/vnd.lucent.voice' }
        .application_vnd_lotus_wordpro { 'application/vnd.lotus-wordpro' }
        .application_x_msmediaview { 'application/x-msmediaview' }
        .video_mpeg { 'video/mpeg' }
        .audio_mpeg { 'audio/mpeg' }
        .audio_x_mpegurl { 'audio/x-mpegurl' }
        .video_vnd_mpegurl { 'video/vnd.mpegurl' }
        .video_x_m4v { 'video/x-m4v' }
        .application_mathematica { 'application/mathematica' }
        .application_vnd_ecowin_chart { 'application/vnd.ecowin.chart' }
        .text_troff { 'text/troff' }
        .application_mathml_xml { 'application/mathml+xml' }
        .text_mathml { 'text/mathml' }
        .application_vnd_sqlite3 { 'application/vnd.sqlite3' }
        .application_vnd_mobius_mbk { 'application/vnd.mobius.mbk' }
        .application_mbox { 'application/mbox' }
        .application_vnd_medcalcdata { 'application/vnd.medcalcdata' }
        .application_vnd_mcd { 'application/vnd.mcd' }
        .text_vnd_curl_mcurl { 'text/vnd.curl.mcurl' }
        .application_x_msaccess { 'application/x-msaccess' }
        .image_vnd_ms_modi { 'image/vnd.ms-modi' }
        .model_mesh { 'model/mesh' }
        .application_vnd_mfmp { 'application/vnd.mfmp' }
        .application_vnd_proteus_magazine { 'application/vnd.proteus.magazine' }
        .application_vnd_mif { 'application/vnd.mif' }
        .video_mj2 { 'video/mj2' }
        .application_vnd_dolby_mlp { 'application/vnd.dolby.mlp' }
        .application_vnd_chipnuts_karaoke_mmd { 'application/vnd.chipnuts.karaoke-mmd' }
        .application_vnd_smaf { 'application/vnd.smaf' }
        .image_vnd_fujixerox_edmics_mmr { 'image/vnd.fujixerox.edmics-mmr' }
        .application_x_msmoney { 'application/x-msmoney' }
        .application_x_mobipocket_ebook { 'application/x-mobipocket-ebook' }
        .video_quicktime { 'video/quicktime' }
        .video_x_sgi_movie { 'video/x-sgi-movie' }
        .video_mp4 { 'video/mp4' }
        .application_x_iso9660_image { 'application/x-iso9660-image' }
        .application_yaml { 'application/yaml' }
        .application_mp4 { 'application/mp4' }
        .application_vnd_mophun_certificate { 'application/vnd.mophun.certificate' }
        .application_vnd_apple_installer_xml { 'application/vnd.apple.installer+xml' }
        .application_vnd_blueice_multipass { 'application/vnd.blueice.multipass' }
        .application_vnd_mophun_application { 'application/vnd.mophun.application' }
        .application_vnd_ms_project { 'application/vnd.ms-project' }
        .application_vnd_ibm_minipay { 'application/vnd.ibm.minipay' }
        .application_vnd_mobius_mqy { 'application/vnd.mobius.mqy' }
        .application_marc { 'application/marc' }
        .application_mediaservercontrol_xml { 'application/mediaservercontrol+xml' }
        .application_vnd_fdsn_mseed { 'application/vnd.fdsn.mseed' }
        .application_vnd_mseq { 'application/vnd.mseq' }
        .application_vnd_epson_msf { 'application/vnd.epson.msf' }
        .application_vnd_mobius_msl { 'application/vnd.mobius.msl' }
        .application_vnd_muvee_style { 'application/vnd.muvee.style' }
        .model_vnd_mts { 'model/vnd.mts' }
        .application_vnd_musician { 'application/vnd.musician' }
        .application_vnd_recordare_musicxml_xml { 'application/vnd.recordare.musicxml+xml' }
        .application_vnd_mfer { 'application/vnd.mfer' }
        .application_mxf { 'application/mxf' }
        .application_vnd_recordare_musicxml { 'application/vnd.recordare.musicxml' }
        .application_xv_xml { 'application/xv+xml' }
        .application_vnd_triscape_mxs { 'application/vnd.triscape.mxs' }
        .application_vnd_nokia_n_gage_symbian_install { 'application/vnd.nokia.n-gage.symbian.install' }
        .application_x_dtbncx_xml { 'application/x-dtbncx+xml' }
        .application_vnd_nokia_n_gage_data { 'application/vnd.nokia.n-gage.data' }
        .application_vnd_neurolanguage_nlu { 'application/vnd.neurolanguage.nlu' }
        .application_vnd_enliven { 'application/vnd.enliven' }
        .application_vnd_noblenet_directory { 'application/vnd.noblenet-directory' }
        .application_vnd_noblenet_sealer { 'application/vnd.noblenet-sealer' }
        .application_vnd_noblenet_web { 'application/vnd.noblenet-web' }
        .image_vnd_net_fpx { 'image/vnd.net-fpx' }
        .application_vnd_lotus_notes { 'application/vnd.lotus-notes' }
        .application_vnd_fujitsu_oasys2 { 'application/vnd.fujitsu.oasys2' }
        .application_vnd_fujitsu_oasys3 { 'application/vnd.fujitsu.oasys3' }
        .application_vnd_fujitsu_oasys { 'application/vnd.fujitsu.oasys' }
        .application_x_msbinder { 'application/x-msbinder' }
        .application_oda { 'application/oda' }
        .application_vnd_oasis_opendocument_database { 'application/vnd.oasis.opendocument.database' }
        .application_vnd_oasis_opendocument_chart { 'application/vnd.oasis.opendocument.chart' }
        .application_vnd_oasis_opendocument_formula { 'application/vnd.oasis.opendocument.formula' }
        .application_vnd_oasis_opendocument_formula_template { 'application/vnd.oasis.opendocument.formula-template' }
        .application_vnd_oasis_opendocument_graphics { 'application/vnd.oasis.opendocument.graphics' }
        .application_vnd_oasis_opendocument_image { 'application/vnd.oasis.opendocument.image' }
        .application_vnd_oasis_opendocument_presentation { 'application/vnd.oasis.opendocument.presentation' }
        .application_vnd_oasis_opendocument_spreadsheet { 'application/vnd.oasis.opendocument.spreadsheet' }
        .application_vnd_oasis_opendocument_text { 'application/vnd.oasis.opendocument.text' }
        .audio_ogg { 'audio/ogg' }
        .video_x_matroska { 'video/x-matroska' }
        .audio_x_matroska { 'audio/x-matroska' }
        .video_ogg { 'video/ogg' }
        .application_ogg { 'application/ogg' }
        .application_onenote { 'application/onenote' }
        .application_oebps_package_xml { 'application/oebps-package+xml' }
        .application_vnd_palm { 'application/vnd.palm' }
        .application_vnd_lotus_organizer { 'application/vnd.lotus-organizer' }
        .application_vnd_yamaha_openscoreformat { 'application/vnd.yamaha.openscoreformat' }
        .application_vnd_yamaha_openscoreformat_osfpvg_xml { 'application/vnd.yamaha.openscoreformat.osfpvg+xml' }
        .application_vnd_oasis_opendocument_chart_template { 'application/vnd.oasis.opendocument.chart-template' }
        .font_woff { 'font/woff' }
        .font_woff2 { 'font/woff2' }
        .application_x_redhat_package_manager { 'application/x-redhat-package-manager' }
        .application_x_perl { 'application/x-perl' }
        .audio_webm { 'audio/webm' }
        .video_webm { 'video/webm' }
        .image_webp { 'image/webp' }
        .application_x_font_otf { 'application/x-font-otf' }
        .font_otf { 'font/otf' }
        .application_vnd_oasis_opendocument_graphics_template { 'application/vnd.oasis.opendocument.graphics-template' }
        .application_vnd_oasis_opendocument_text_web { 'application/vnd.oasis.opendocument.text-web' }
        .application_vnd_oasis_opendocument_image_template { 'application/vnd.oasis.opendocument.image-template' }
        .application_vnd_oasis_opendocument_text_master { 'application/vnd.oasis.opendocument.text-master' }
        .application_vnd_oasis_opendocument_presentation_template { 'application/vnd.oasis.opendocument.presentation-template' }
        .application_vnd_oasis_opendocument_spreadsheet_template { 'application/vnd.oasis.opendocument.spreadsheet-template' }
        .application_vnd_oasis_opendocument_text_template { 'application/vnd.oasis.opendocument.text-template' }
        .application_vnd_openofficeorg_extension { 'application/vnd.openofficeorg.extension' }
        .text_x_pascal { 'text/x-pascal' }
        .application_pkcs10 { 'application/pkcs10' }
        .application_x_pkcs12 { 'application/x-pkcs12' }
        .application_x_pkcs7_certificates { 'application/x-pkcs7-certificates' }
        .application_pkcs7_mime { 'application/pkcs7-mime' }
        .application_x_pkcs7_certreqresp { 'application/x-pkcs7-certreqresp' }
        .application_pkcs7_signature { 'application/pkcs7-signature' }
        .application_vnd_powerbuilder6 { 'application/vnd.powerbuilder6' }
        .image_x_portable_bitmap { 'image/x-portable-bitmap' }
        .application_x_font_pcf { 'application/x-font-pcf' }
        .application_vnd_hp_pcl { 'application/vnd.hp-pcl' }
        .application_vnd_hp_pclxl { 'application/vnd.hp-pclxl' }
        .image_x_pict { 'image/x-pict' }
        .application_vnd_curl_pcurl { 'application/vnd.curl.pcurl' }
        .image_x_pcx { 'image/x-pcx' }
        .application_pdf { 'application/pdf' }
        .application_font_tdpfr { 'application/font-tdpfr' }
        .image_x_portable_graymap { 'image/x-portable-graymap' }
        .application_x_chess_pgn { 'application/x-chess-pgn' }
        .application_pgp_encrypted { 'application/pgp-encrypted' }
        .application_pkixcmp { 'application/pkixcmp' }
        .application_pkix_pkipath { 'application/pkix-pkipath' }
        .application_vnd_3gpp_pic_bw_large { 'application/vnd.3gpp.pic-bw-large' }
        .application_vnd_mobius_plc { 'application/vnd.mobius.plc' }
        .application_vnd_pocketlearn { 'application/vnd.pocketlearn' }
        .application_pls_xml { 'application/pls+xml' }
        .application_vnd_ctc_posml { 'application/vnd.ctc-posml' }
        .image_png { 'image/png' }
        .image_x_portable_anymap { 'image/x-portable-anymap' }
        .application_vnd_macports_portpkg { 'application/vnd.macports.portpkg' }
        .application_vnd_ms_powerpoint { 'application/vnd.ms-powerpoint' }
        .application_vnd_ms_powerpoint_template_macroenabled_12 { 'application/vnd.ms-powerpoint.template.macroenabled.12' }
        .application_vnd_openxmlformats_officedocument_presentationml_template { 'application/vnd.openxmlformats-officedocument.presentationml.template' }
        .application_vnd_ms_powerpoint_addin_macroenabled_12 { 'application/vnd.ms-powerpoint.addin.macroenabled.12' }
        .application_vnd_cups_ppd { 'application/vnd.cups-ppd' }
        .image_x_portable_pixmap { 'image/x-portable-pixmap' }
        .application_vnd_ms_powerpoint_slideshow_macroenabled_12 { 'application/vnd.ms-powerpoint.slideshow.macroenabled.12' }
        .application_vnd_openxmlformats_officedocument_presentationml_slideshow { 'application/vnd.openxmlformats-officedocument.presentationml.slideshow' }
        .application_vnd_ms_powerpoint_presentation_macroenabled_12 { 'application/vnd.ms-powerpoint.presentation.macroenabled.12' }
        .application_vnd_openxmlformats_officedocument_presentationml_presentation { 'application/vnd.openxmlformats-officedocument.presentationml.presentation' }
        .application_vnd_lotus_freelance { 'application/vnd.lotus-freelance' }
        .application_pics_rules { 'application/pics-rules' }
        .application_prql { 'application/prql' }
        .application_vnd_3gpp_pic_bw_small { 'application/vnd.3gpp.pic-bw-small' }
        .image_vnd_adobe_photoshop { 'image/vnd.adobe.photoshop' }
        .application_x_font_linux_psf { 'application/x-font-linux-psf' }
        .application_vnd_pvi_ptid1 { 'application/vnd.pvi.ptid1' }
        .application_x_mspublisher { 'application/x-mspublisher' }
        .application_vnd_3gpp_pic_bw_var { 'application/vnd.3gpp.pic-bw-var' }
        .application_vnd_3m_post_it_notes { 'application/vnd.3m.post-it-notes' }
        .text_x_python { 'text/x-python' }
        .audio_vnd_ms_playready_media_pya { 'audio/vnd.ms-playready.media.pya' }
        .video_vnd_ms_playready_media_pyv { 'video/vnd.ms-playready.media.pyv' }
        .application_vnd_epson_quickanime { 'application/vnd.epson.quickanime' }
        .application_vnd_intu_qbo { 'application/vnd.intu.qbo' }
        .application_vnd_intu_qfx { 'application/vnd.intu.qfx' }
        .application_vnd_publishare_delta_tree { 'application/vnd.publishare-delta-tree' }
        .application_vnd_quark_quarkxpress { 'application/vnd.quark.quarkxpress' }
        .audio_x_pn_realaudio { 'audio/x-pn-realaudio' }
        .application_vnd_rar { 'application/vnd.rar' }
        .application_x_rar_compressed { 'application/x-rar-compressed' }
        .image_x_cmu_raster { 'image/x-cmu-raster' }
        .application_vnd_ipunplugged_rcprofile { 'application/vnd.ipunplugged.rcprofile' }
        .application_rdf_xml { 'application/rdf+xml' }
        .application_vnd_data_vision_rdz { 'application/vnd.data-vision.rdz' }
        .application_vnd_businessobjects { 'application/vnd.businessobjects' }
        .application_x_dtbresource_xml { 'application/x-dtbresource+xml' }
        .image_x_rgb { 'image/x-rgb' }
        .application_reginfo_xml { 'application/reginfo+xml' }
        .application_resource_lists_xml { 'application/resource-lists+xml' }
        .image_vnd_fujixerox_edmics_rlc { 'image/vnd.fujixerox.edmics-rlc' }
        .application_resource_lists_diff_xml { 'application/resource-lists-diff+xml' }
        .application_vnd_rn_realmedia { 'application/vnd.rn-realmedia' }
        .audio_x_pn_realaudio_plugin { 'audio/x-pn-realaudio-plugin' }
        .application_vnd_jcp_javame_midlet_rms { 'application/vnd.jcp.javame.midlet-rms' }
        .application_relax_ng_compact_syntax { 'application/relax-ng-compact-syntax' }
        .application_x_rpm { 'application/x-rpm' }
        .application_vnd_nokia_radio_presets { 'application/vnd.nokia.radio-presets' }
        .application_vnd_nokia_radio_preset { 'application/vnd.nokia.radio-preset' }
        .application_sparql_query { 'application/sparql-query' }
        .application_rls_services_xml { 'application/rls-services+xml' }
        .application_rsd_xml { 'application/rsd+xml' }
        .application_rss_xml { 'application/rss+xml' }
        .application_rtf { 'application/rtf' }
        .text_richtext { 'text/richtext' }
        .application_vnd_yamaha_smaf_audio { 'application/vnd.yamaha.smaf-audio' }
        .application_sbml_xml { 'application/sbml+xml' }
        .application_vnd_ibm_secure_container { 'application/vnd.ibm.secure-container' }
        .application_x_msschedule { 'application/x-msschedule' }
        .application_vnd_lotus_screencam { 'application/vnd.lotus-screencam' }
        .application_scvp_cv_request { 'application/scvp-cv-request' }
        .application_scvp_cv_response { 'application/scvp-cv-response' }
        .text_vnd_curl_scurl { 'text/vnd.curl.scurl' }
        .application_vnd_stardivision_draw { 'application/vnd.stardivision.draw' }
        .application_vnd_stardivision_calc { 'application/vnd.stardivision.calc' }
        .application_vnd_stardivision_impress { 'application/vnd.stardivision.impress' }
        .application_vnd_solent_sdkm_xml { 'application/vnd.solent.sdkm+xml' }
        .application_sdp { 'application/sdp' }
        .application_vnd_stardivision_writer { 'application/vnd.stardivision.writer' }
        .application_vnd_seemail { 'application/vnd.seemail' }
        .application_vnd_sema { 'application/vnd.sema' }
        .application_vnd_semd { 'application/vnd.semd' }
        .application_vnd_semf { 'application/vnd.semf' }
        .application_java_serialized_object { 'application/java-serialized-object' }
        .application_set_payment_initiation { 'application/set-payment-initiation' }
        .application_set_registration_initiation { 'application/set-registration-initiation' }
        .application_vnd_hydrostatix_sof_data { 'application/vnd.hydrostatix.sof-data' }
        .application_vnd_spotfire_sfs { 'application/vnd.spotfire.sfs' }
        .application_vnd_stardivision_writer_global { 'application/vnd.stardivision.writer-global' }
        .text_sgml { 'text/sgml' }
        .application_x_sh { 'application/x-sh' }
        .application_x_shar { 'application/x-shar' }
        .application_shf_xml { 'application/shf+xml' }
        .text_vnd_wap_si { 'text/vnd.wap.si' }
        .application_vnd_wap_sic { 'application/vnd.wap.sic' }
        .application_vnd_symbian_install { 'application/vnd.symbian.install' }
        .application_x_stuffit { 'application/x-stuffit' }
        .application_x_stuffitx { 'application/x-stuffitx' }
        .application_vnd_koan { 'application/vnd.koan' }
        .text_vnd_wap_sl { 'text/vnd.wap.sl' }
        .application_vnd_wap_slc { 'application/vnd.wap.slc' }
        .application_vnd_ms_powerpoint_slide_macroenabled_12 { 'application/vnd.ms-powerpoint.slide.macroenabled.12' }
        .application_vnd_openxmlformats_officedocument_presentationml_slide { 'application/vnd.openxmlformats-officedocument.presentationml.slide' }
        .application_vnd_epson_salt { 'application/vnd.epson.salt' }
        .application_vnd_stardivision_math { 'application/vnd.stardivision.math' }
        .application_smil_xml { 'application/smil+xml' }
        .application_x_font_snf { 'application/x-font-snf' }
        .application_vnd_yamaha_smaf_phrase { 'application/vnd.yamaha.smaf-phrase' }
        .application_x_futuresplash { 'application/x-futuresplash' }
        .text_vnd_in3d_spot { 'text/vnd.in3d.spot' }
        .application_scvp_vp_response { 'application/scvp-vp-response' }
        .application_scvp_vp_request { 'application/scvp-vp-request' }
        .application_x_wais_source { 'application/x-wais-source' }
        .application_sparql_results_xml { 'application/sparql-results+xml' }
        .application_vnd_kodak_descriptor { 'application/vnd.kodak-descriptor' }
        .application_vnd_epson_ssf { 'application/vnd.epson.ssf' }
        .application_ssml_xml { 'application/ssml+xml' }
        .application_vnd_sun_xml_calc_template { 'application/vnd.sun.xml.calc.template' }
        .application_vnd_sun_xml_draw_template { 'application/vnd.sun.xml.draw.template' }
        .application_vnd_wt_stf { 'application/vnd.wt.stf' }
        .application_vnd_sun_xml_impress_template { 'application/vnd.sun.xml.impress.template' }
        .application_hyperstudio { 'application/hyperstudio' }
        .application_vnd_ms_pki_stl { 'application/vnd.ms-pki.stl' }
        .application_vnd_pg_format { 'application/vnd.pg.format' }
        .application_vnd_sun_xml_writer_template { 'application/vnd.sun.xml.writer.template' }
        .application_vnd_sus_calendar { 'application/vnd.sus-calendar' }
        .application_x_sv4cpio { 'application/x-sv4cpio' }
        .application_x_sv4crc { 'application/x-sv4crc' }
        .application_vnd_svd { 'application/vnd.svd' }
        .image_svg_xml { 'image/svg+xml' }
        .application_x_shockwave_flash { 'application/x-shockwave-flash' }
        .application_vnd_arastra_swi { 'application/vnd.arastra.swi' }
        .application_vnd_sun_xml_calc { 'application/vnd.sun.xml.calc' }
        .application_vnd_sun_xml_draw { 'application/vnd.sun.xml.draw' }
        .application_vnd_sun_xml_writer_global { 'application/vnd.sun.xml.writer.global' }
        .application_vnd_sun_xml_impress { 'application/vnd.sun.xml.impress' }
        .application_vnd_sun_xml_math { 'application/vnd.sun.xml.math' }
        .application_vnd_sun_xml_writer { 'application/vnd.sun.xml.writer' }
        .application_vnd_tao_intent_module_archive { 'application/vnd.tao.intent-module-archive' }
        .application_x_tar { 'application/x-tar' }
        .application_vnd_3gpp2_tcap { 'application/vnd.3gpp2.tcap' }
        .application_x_tcl { 'application/x-tcl' }
        .application_vnd_smart_teacher { 'application/vnd.smart.teacher' }
        .application_x_tex { 'application/x-tex' }
        .application_x_texinfo { 'application/x-texinfo' }
        .application_x_tex_tfm { 'application/x-tex-tfm' }
        .image_tiff { 'image/tiff' }
        .application_vnd_tmobile_livetv { 'application/vnd.tmobile-livetv' }
        .application_x_bittorrent { 'application/x-bittorrent' }
        .application_vnd_groove_tool_template { 'application/vnd.groove-tool-template' }
        .application_vnd_trid_tpt { 'application/vnd.trid.tpt' }
        .application_vnd_trueapp { 'application/vnd.trueapp' }
        .application_x_msterminal { 'application/x-msterminal' }
        .text_tab_separated_values { 'text/tab-separated-values' }
        .application_x_font_ttf { 'application/x-font-ttf' }
        .application_vnd_simtech_mindmapper { 'application/vnd.simtech-mindmapper' }
        .application_vnd_genomatix_tuxedo { 'application/vnd.genomatix.tuxedo' }
        .application_vnd_mobius_txf { 'application/vnd.mobius.txf' }
        .application_vnd_ufdl { 'application/vnd.ufdl' }
        .test_mimetype { 'test/mimetype' }
        .application_vnd_umajin { 'application/vnd.umajin' }
        .application_vnd_unity { 'application/vnd.unity' }
        .application_vnd_uoml_xml { 'application/vnd.uoml+xml' }
        .text_uri_list { 'text/uri-list' }
        .application_x_ustar { 'application/x-ustar' }
        .application_vnd_uiq_theme { 'application/vnd.uiq.theme' }
        .text_x_uuencode { 'text/x-uuencode' }
        .application_x_cdlink { 'application/x-cdlink' }
        .text_x_vcard { 'text/x-vcard' }
        .application_vnd_groove_vcard { 'application/vnd.groove-vcard' }
        .text_x_vcalendar { 'text/x-vcalendar' }
        .application_vnd_vcx { 'application/vnd.vcx' }
        .application_vnd_visionary { 'application/vnd.visionary' }
        .video_vnd_vivo { 'video/vnd.vivo' }
        .model_vrml { 'model/vrml' }
        .application_vnd_visio { 'application/vnd.visio' }
        .application_vnd_vsf { 'application/vnd.vsf' }
        .model_vnd_vtu { 'model/vnd.vtu' }
        .application_voicexml_xml { 'application/voicexml+xml' }
        .application_x_doom { 'application/x-doom' }
        .video_mp2t { 'video/mp2t' }
        .audio_vnd_wav { 'audio/vnd.wav' }
        .audio_x_ms_wax { 'audio/x-ms-wax' }
        .image_vnd_wap_wbmp { 'image/vnd.wap.wbmp' }
        .application_vnd_criticaltools_wbs_xml { 'application/vnd.criticaltools.wbs+xml' }
        .application_vnd_wap_wbxml { 'application/vnd.wap.wbxml' }
        .application_vnd_ms_works { 'application/vnd.ms-works' }
        .video_x_ms_wm { 'video/x-ms-wm' }
        .audio_x_ms_wma { 'audio/x-ms-wma' }
        .application_x_ms_wmd { 'application/x-ms-wmd' }
        .application_x_msmetafile { 'application/x-msmetafile' }
        .text_vnd_wap_wml { 'text/vnd.wap.wml' }
        .application_vnd_wap_wmlc { 'application/vnd.wap.wmlc' }
        .text_vnd_wap_wmlscript { 'text/vnd.wap.wmlscript' }
        .application_vnd_wap_wmlscriptc { 'application/vnd.wap.wmlscriptc' }
        .video_x_ms_wmv { 'video/x-ms-wmv' }
        .video_x_ms_wmx { 'video/x-ms-wmx' }
        .application_x_ms_wmz { 'application/x-ms-wmz' }
        .application_vnd_wordperfect { 'application/vnd.wordperfect' }
        .application_vnd_ms_wpl { 'application/vnd.ms-wpl' }
        .application_vnd_wqd { 'application/vnd.wqd' }
        .application_x_mswrite { 'application/x-mswrite' }
        .application_wsdl_xml { 'application/wsdl+xml' }
        .application_wspolicy_xml { 'application/wspolicy+xml' }
        .application_vnd_webturbo { 'application/vnd.webturbo' }
        .video_x_ms_wvx { 'video/x-ms-wvx' }
        .application_vnd_hzn_3d_crossword { 'application/vnd.hzn-3d-crossword' }
        .application_x_silverlight_app { 'application/x-silverlight-app' }
        .application_vnd_xara { 'application/vnd.xara' }
        .application_x_ms_xbap { 'application/x-ms-xbap' }
        .application_vnd_fujixerox_docuworks_binder { 'application/vnd.fujixerox.docuworks.binder' }
        .image_x_xbitmap { 'image/x-xbitmap' }
        .application_vnd_syncml_dm_xml { 'application/vnd.syncml.dm+xml' }
        .application_vnd_adobe_xdp_xml { 'application/vnd.adobe.xdp+xml' }
        .application_vnd_fujixerox_docuworks { 'application/vnd.fujixerox.docuworks' }
        .application_xenc_xml { 'application/xenc+xml' }
        .application_patch_ops_error_xml { 'application/patch-ops-error+xml' }
        .application_vnd_adobe_xfdf { 'application/vnd.adobe.xfdf' }
        .application_vnd_xfdl { 'application/vnd.xfdl' }
        .application_xhtml_xml { 'application/xhtml+xml' }
        .image_vnd_xiff { 'image/vnd.xiff' }
        .application_vnd_ms_excel { 'application/vnd.ms-excel' }
        .application_vnd_ms_excel_addin_macroenabled_12 { 'application/vnd.ms-excel.addin.macroenabled.12' }
        .application_vnd_ms_excel_sheet_binary_macroenabled_12 { 'application/vnd.ms-excel.sheet.binary.macroenabled.12' }
        .application_vnd_ms_excel_sheet_macroenabled_12 { 'application/vnd.ms-excel.sheet.macroenabled.12' }
        .application_vnd_openxmlformats_officedocument_spreadsheetml_sheet { 'application/vnd.openxmlformats-officedocument.spreadsheetml.sheet' }
        .application_vnd_ms_excel_template_macroenabled_12 { 'application/vnd.ms-excel.template.macroenabled.12' }
        .application_vnd_openxmlformats_officedocument_spreadsheetml_template { 'application/vnd.openxmlformats-officedocument.spreadsheetml.template' }
        .application_xml { 'application/xml' }
        .application_vnd_olpc_sugar { 'application/vnd.olpc-sugar' }
        .application_xop_xml { 'application/xop+xml' }
        .application_x_xpinstall { 'application/x-xpinstall' }
        .image_x_xpixmap { 'image/x-xpixmap' }
        .application_vnd_is_xpr { 'application/vnd.is-xpr' }
        .application_vnd_ms_xpsdocument { 'application/vnd.ms-xpsdocument' }
        .application_vnd_intercon_formnet { 'application/vnd.intercon.formnet' }
        .application_xslt_xml { 'application/xslt+xml' }
        .application_vnd_syncml_xml { 'application/vnd.syncml+xml' }
        .application_xspf_xml { 'application/xspf+xml' }
        .application_vnd_mozilla_xul_xml { 'application/vnd.mozilla.xul+xml' }
        .image_x_xwindowdump { 'image/x-xwindowdump' }
        .chemical_x_xyz { 'chemical/x-xyz' }
        .application_vnd_zzazz_deck_xml { 'application/vnd.zzazz.deck+xml' }
        .application_zip { 'application/zip' }
        .application_x_zip_compressed { 'application/x-zip-compressed' }
        .application_zip_compressed { 'application/zip-compressed' }
        .application_vnd_zul { 'application/vnd.zul' }
        .application_vnd_handheld_entertainment_xml { 'application/vnd.handheld-entertainment+xml' }
        .image_x_adobe_dng { 'image/x-adobe-dng' }
        .image_x_sony_arw { 'image/x-sony-arw' }
        .image_x_canon_cr2 { 'image/x-canon-cr2' }
        .image_x_canon_crw { 'image/x-canon-crw' }
        .image_x_kodak_dcr { 'image/x-kodak-dcr' }
        .image_x_epson_erf { 'image/x-epson-erf' }
        .image_x_kodak_k25 { 'image/x-kodak-k25' }
        .image_x_kodak_kdc { 'image/x-kodak-kdc' }
        .image_x_minolta_mrw { 'image/x-minolta-mrw' }
        .image_x_nikon_nef { 'image/x-nikon-nef' }
        .image_x_olympus_orf { 'image/x-olympus-orf' }
        .image_x_pentax_pef { 'image/x-pentax-pef' }
        .image_x_fuji_raf { 'image/x-fuji-raf' }
        .image_x_panasonic_raw { 'image/x-panasonic-raw' }
        .audio_flac { 'audio/flac' }
        .image_x_sony_sr2 { 'image/x-sony-sr2' }
        .image_x_sony_srf { 'image/x-sony-srf' }
        .image_x_sigma_x3f { 'image/x-sigma-x3f' }
    }
}
