module mime

pub fn Mime.from_extension(extension string) ?Mime {
    return match extension {
        '123' { Mime.application_vnd_lotus_1_2_3 }
        '3dml' { Mime.text_vnd_in3d_3dml }
        '3g2' { Mime.video_3gpp2 }
        '3ga' { Mime.audio_mp4 }
        '3gp' { Mime.video_3gpp }
        '3gp2' { Mime.audio_mp4 }
        '3gpa' { Mime.audio_mp4 }
        '3gpp' { Mime.audio_mp4 }
        '3gpp2' { Mime.audio_mp4 }
        '7z' { Mime.application_x_7z_compressed }
        'a' { Mime.application_octet_stream }
        'aab' { Mime.application_x_authorware_bin }
        'aac' { Mime.audio_aac }
        'aacp' { Mime.audio_aacp }
        'aam' { Mime.application_x_authorware_map }
        'aas' { Mime.application_x_authorware_seg }
        'abw' { Mime.application_x_abiword }
        'abw.gz' { Mime.application_x_abiword }
        'acc' { Mime.application_vnd_americandynamics_acc }
        'ace' { Mime.application_x_ace_compressed }
        'acu' { Mime.application_vnd_acucobol }
        'acutc' { Mime.application_vnd_acucorp }
        'adp' { Mime.audio_adpcm }
        'aep' { Mime.application_vnd_audiograph }
        'aff' { Mime.audio_aiff }
        'afm' { Mime.application_x_font_type1 }
        'afp' { Mime.application_vnd_ibm_modcap }
        'ai' { Mime.application_postscript }
        'aif' { Mime.audio_aiff }
        'aiff' { Mime.audio_aiff }
        'air' { Mime.application_vnd_adobe_air_application_installer_package_zip }
        'ami' { Mime.application_vnd_amiga_ami }
        'apk' { Mime.application_vnd_android_package_archive }
        'application' { Mime.application_x_ms_application }
        'apr' { Mime.application_vnd_lotus_approach }
        'arw' { Mime.image_x_sony_arw }
        'asc' { Mime.application_pgp_signature }
        'asf' { Mime.video_x_ms_asf }
        'asm' { Mime.text_x_asm }
        'aso' { Mime.application_vnd_accpac_simply_aso }
        'asx' { Mime.video_x_ms_asf }
        'atc' { Mime.application_vnd_acucorp }
        'atom' { Mime.application_atom_xml }
        'atomcat' { Mime.application_atomcat_xml }
        'atomsvc' { Mime.application_atomsvc_xml }
        'atx' { Mime.application_vnd_antix_game_component }
        'au' { Mime.audio_basic }
        'avi' { Mime.video_x_msvideo }
        'avif' { Mime.image_avif }
        'avifs' { Mime.image_avif_sequence }
        'aw' { Mime.application_applixware }
        'azf' { Mime.application_vnd_airzip_filesecure_azf }
        'azs' { Mime.application_vnd_airzip_filesecure_azs }
        'azw' { Mime.application_vnd_amazon_ebook }
        'bat' { Mime.application_x_msdownload }
        'bcpio' { Mime.application_x_bcpio }
        'bdf' { Mime.application_x_font_bdf }
        'bdm' { Mime.application_vnd_syncml_dm_wbxml }
        'bh2' { Mime.application_vnd_fujitsu_oasysprs }
        'bin' { Mime.application_octet_stream }
        'bmi' { Mime.application_vnd_bmi }
        'bmp' { Mime.image_bmp }
        'book' { Mime.application_vnd_framemaker }
        'box' { Mime.application_vnd_previewsystems_box }
        'boz' { Mime.application_x_bzip2 }
        'bpk' { Mime.application_octet_stream }
        'btif' { Mime.image_prs_btif }
        'bz' { Mime.application_x_bzip }
        'bz2' { Mime.application_x_bzip2 }
        'c' { Mime.text_x_c }
        'c4d' { Mime.application_vnd_clonk_c4group }
        'c4f' { Mime.application_vnd_clonk_c4group }
        'c4g' { Mime.application_vnd_clonk_c4group }
        'c4p' { Mime.application_vnd_clonk_c4group }
        'c4u' { Mime.application_vnd_clonk_c4group }
        'cab' { Mime.application_vnd_ms_cab_compressed }
        'car' { Mime.application_vnd_curl_car }
        'cat' { Mime.application_vnd_ms_pki_seccat }
        'cc' { Mime.text_x_c }
        'cct' { Mime.application_x_director }
        'ccxml' { Mime.application_ccxml_xml }
        'cdbcmsg' { Mime.application_vnd_contact_cmsg }
        'cdf' { Mime.application_x_netcdf }
        'cdkey' { Mime.application_vnd_mediastation_cdkey }
        'cdr' { Mime.application_x_iso9660_image }
        'cdx' { Mime.chemical_x_cdx }
        'cdxml' { Mime.application_vnd_chemdraw_xml }
        'cdy' { Mime.application_vnd_cinderella }
        'cer' { Mime.application_pkix_cert }
        'cgm' { Mime.image_cgm }
        'chat' { Mime.application_x_chat }
        'chm' { Mime.application_vnd_ms_htmlhelp }
        'chrt' { Mime.application_vnd_kde_kchart }
        'cif' { Mime.chemical_x_cif }
        'cii' { Mime.application_vnd_anser_web_certificate_issue_initiation }
        'cil' { Mime.application_vnd_ms_artgalry }
        'cla' { Mime.application_vnd_claymore }
        'class' { Mime.application_java_vm }
        'clkk' { Mime.application_vnd_crick_clicker_keyboard }
        'clkp' { Mime.application_vnd_crick_clicker_palette }
        'clkt' { Mime.application_vnd_crick_clicker_template }
        'clkw' { Mime.application_vnd_crick_clicker_wordbank }
        'clkx' { Mime.application_vnd_crick_clicker }
        'clp' { Mime.application_x_msclip }
        'cmc' { Mime.application_vnd_cosmocaller }
        'cmdf' { Mime.chemical_x_cmdf }
        'cml' { Mime.chemical_x_cml }
        'cmp' { Mime.application_vnd_yellowriver_custom_menu }
        'cmx' { Mime.image_x_cmx }
        'cod' { Mime.application_vnd_rim_cod }
        'com' { Mime.application_x_msdownload }
        'conf' { Mime.text_plain }
        'cpio' { Mime.application_x_cpio }
        'cpp' { Mime.text_x_c }
        'cpt' { Mime.application_mac_compactpro }
        'cr2' { Mime.image_x_canon_cr2 }
        'crd' { Mime.application_x_mscardfile }
        'crl' { Mime.application_pkix_crl }
        'crt' { Mime.application_x_x509_ca_cert }
        'crw' { Mime.image_x_canon_crw }
        'csh' { Mime.application_x_csh }
        'csml' { Mime.chemical_x_csml }
        'csp' { Mime.application_vnd_commonspace }
        'css' { Mime.text_css }
        'cst' { Mime.application_x_director }
        'csv' { Mime.text_csv }
        'cu' { Mime.application_cu_seeme }
        'curl' { Mime.text_vnd_curl }
        'cww' { Mime.application_prs_cww }
        'cxt' { Mime.application_x_director }
        'cxx' { Mime.text_x_c }
        'daf' { Mime.application_vnd_mobius_daf }
        'dataless' { Mime.application_vnd_fdsn_seed }
        'davmount' { Mime.application_davmount_xml }
        'db' { Mime.application_vnd_sqlite3 }
        'db-shm' { Mime.application_vnd_sqlite3 }
        'db-wal' { Mime.application_vnd_sqlite3 }
        'dcr' { Mime.application_x_director }
        'dcurl' { Mime.text_vnd_curl_dcurl }
        'dd2' { Mime.application_vnd_oma_dd2_xml }
        'ddd' { Mime.application_vnd_fujixerox_ddd }
        'deb' { Mime.application_vnd_debian_binary_package }
        'def' { Mime.text_plain }
        'deploy' { Mime.application_octet_stream }
        'der' { Mime.application_x_x509_ca_cert }
        'dfac' { Mime.application_vnd_dreamfactory }
        'dic' { Mime.text_x_c }
        'diff' { Mime.text_plain }
        'dir' { Mime.application_x_director }
        'dis' { Mime.application_vnd_mobius_dis }
        'dist' { Mime.application_octet_stream }
        'distz' { Mime.application_octet_stream }
        'djv' { Mime.image_vnd_djvu }
        'djvu' { Mime.image_vnd_djvu }
        'dll' { Mime.application_x_msdownload }
        'dmg' { Mime.application_octet_stream }
        'dms' { Mime.application_octet_stream }
        'dna' { Mime.application_vnd_dna }
        'dng' { Mime.image_x_adobe_dng }
        'doc' { Mime.application_msword }
        'docm' { Mime.application_vnd_ms_word_document_macroenabled_12 }
        'docx' { Mime.application_vnd_openxmlformats_officedocument_wordprocessingml_document }
        'dot' { Mime.application_msword }
        'dotm' { Mime.application_vnd_ms_word_template_macroenabled_12 }
        'dotx' { Mime.application_vnd_openxmlformats_officedocument_wordprocessingml_template }
        'dp' { Mime.application_vnd_osgi_dp }
        'dpg' { Mime.application_vnd_dpgraph }
        'dsc' { Mime.text_prs_lines_tag }
        'dtb' { Mime.application_x_dtbook_xml }
        'dtd' { Mime.application_xml_dtd }
        'dts' { Mime.audio_vnd_dts }
        'dtshd' { Mime.audio_vnd_dts_hd }
        'dump' { Mime.application_octet_stream }
        'dvi' { Mime.application_x_dvi }
        'dwf' { Mime.model_vnd_dwf }
        'dwg' { Mime.image_vnd_dwg }
        'dxf' { Mime.image_vnd_dxf }
        'dxp' { Mime.application_vnd_spotfire_dxp }
        'dxr' { Mime.application_x_director }
        'ecelp4800' { Mime.audio_vnd_nuera_ecelp4800 }
        'ecelp7470' { Mime.audio_vnd_nuera_ecelp7470 }
        'ecelp9600' { Mime.audio_vnd_nuera_ecelp9600 }
        'ecma' { Mime.application_ecmascript }
        'edm' { Mime.application_vnd_novadigm_edm }
        'edx' { Mime.application_vnd_novadigm_edx }
        'efif' { Mime.application_vnd_picsel }
        'ei6' { Mime.application_vnd_pg_osasli }
        'elc' { Mime.application_octet_stream }
        'eml' { Mime.message_rfc822 }
        'emma' { Mime.application_emma_xml }
        'eol' { Mime.audio_vnd_digital_winds }
        'eot' { Mime.application_vnd_ms_fontobject }
        'eps' { Mime.application_postscript }
        'epub' { Mime.application_epub_zip }
        'erf' { Mime.image_x_epson_erf }
        'es3' { Mime.application_vnd_eszigno3_xml }
        'esf' { Mime.application_vnd_epson_esf }
        'et3' { Mime.application_vnd_eszigno3_xml }
        'etx' { Mime.text_x_setext }
        'exe' { Mime.application_x_msdownload }
        'ext' { Mime.application_vnd_novadigm_ext }
        'ez' { Mime.application_andrew_inset }
        'ez2' { Mime.application_vnd_ezpix_album }
        'ez3' { Mime.application_vnd_ezpix_package }
        'f' { Mime.text_x_fortran }
        'f4v' { Mime.video_x_f4v }
        'f77' { Mime.text_x_fortran }
        'f90' { Mime.text_x_fortran }
        'fbs' { Mime.image_vnd_fastbidsheet }
        'fdf' { Mime.application_vnd_fdf }
        'fe_launch' { Mime.application_vnd_denovo_fcselayout_link }
        'fg5' { Mime.application_vnd_fujitsu_oasysgp }
        'fgd' { Mime.application_x_director }
        'fh' { Mime.image_x_freehand }
        'fh4' { Mime.image_x_freehand }
        'fh5' { Mime.image_x_freehand }
        'fh7' { Mime.image_x_freehand }
        'fhc' { Mime.image_x_freehand }
        'fig' { Mime.application_x_xfig }
        'flac' { Mime.audio_flac }
        'fli' { Mime.video_x_fli }
        'flo' { Mime.application_vnd_micrografx_flo }
        'flv' { Mime.video_x_flv }
        'flw' { Mime.application_vnd_kde_kivio }
        'flx' { Mime.text_vnd_fmi_flexstor }
        'fly' { Mime.text_vnd_fly }
        'fm' { Mime.application_vnd_framemaker }
        'fnc' { Mime.application_vnd_frogans_fnc }
        'for' { Mime.text_x_fortran }
        'fpx' { Mime.image_vnd_fpx }
        'frame' { Mime.application_vnd_framemaker }
        'fsc' { Mime.application_vnd_fsc_weblaunch }
        'fst' { Mime.image_vnd_fst }
        'ftc' { Mime.application_vnd_fluxtime_clip }
        'fti' { Mime.application_vnd_anser_web_funds_transfer_initiation }
        'fvt' { Mime.video_vnd_fvt }
        'fzs' { Mime.application_vnd_fuzzysheet }
        'g3' { Mime.image_g3fax }
        'gac' { Mime.application_vnd_groove_account }
        'gbr' { Mime.application_vnd_gerber }
        'gcode' { Mime.gcode }
        'gdl' { Mime.model_vnd_gdl }
        'geo' { Mime.application_vnd_dynageo }
        'gex' { Mime.application_vnd_geometry_explorer }
        'ggb' { Mime.application_vnd_geogebra_file }
        'ggt' { Mime.application_vnd_geogebra_tool }
        'ghf' { Mime.application_vnd_groove_help }
        'gif' { Mime.image_gif }
        'gim' { Mime.application_vnd_groove_identity_message }
        'gmx' { Mime.application_vnd_gmx }
        'gnumeric' { Mime.application_x_gnumeric }
        'gph' { Mime.application_vnd_flographit }
        'gqf' { Mime.application_vnd_grafeq }
        'gqs' { Mime.application_vnd_grafeq }
        'gram' { Mime.application_srgs }
        'gre' { Mime.application_vnd_geometry_explorer }
        'grv' { Mime.application_vnd_groove_injector }
        'grxml' { Mime.application_srgs_xml }
        'gsf' { Mime.application_x_font_ghostscript }
        'gtar' { Mime.application_x_gtar }
        'gtm' { Mime.application_vnd_groove_tool_message }
        'gtw' { Mime.model_vnd_gtw }
        'gv' { Mime.text_vnd_graphviz }
        'gz' { Mime.application_x_gzip }
        'h' { Mime.text_x_c }
        'h261' { Mime.video_h261 }
        'h263' { Mime.video_h263 }
        'h264' { Mime.video_h264 }
        'hbci' { Mime.application_vnd_hbci }
        'hdf' { Mime.application_x_hdf }
        'heic' { Mime.image_heic }
        'heif' { Mime.image_heic }
        'hh' { Mime.text_x_c }
        'hlp' { Mime.application_winhlp }
        'hpgl' { Mime.application_vnd_hp_hpgl }
        'hpid' { Mime.application_vnd_hp_hpid }
        'hps' { Mime.application_vnd_hp_hps }
        'hqx' { Mime.application_mac_binhex40 }
        'htke' { Mime.application_vnd_kenameaapp }
        'htm' { Mime.text_html }
        'html' { Mime.text_html }
        'hvd' { Mime.application_vnd_yamaha_hv_dic }
        'hvp' { Mime.application_vnd_yamaha_hv_voice }
        'hvs' { Mime.application_vnd_yamaha_hv_script }
        'icc' { Mime.application_vnd_iccprofile }
        'ice' { Mime.x_conference_x_cooltalk }
        'icm' { Mime.application_vnd_iccprofile }
        'icns' { Mime.image_x_icns }
        'ico' { Mime.image_x_icon }
        'ics' { Mime.text_calendar }
        'ief' { Mime.image_ief }
        'ifb' { Mime.text_calendar }
        'ifm' { Mime.application_vnd_shana_informed_formdata }
        'iges' { Mime.model_iges }
        'igl' { Mime.application_vnd_igloader }
        'igs' { Mime.model_iges }
        'igx' { Mime.application_vnd_micrografx_igx }
        'iif' { Mime.application_vnd_shana_informed_interchange }
        'imp' { Mime.application_vnd_accpac_simply_imp }
        'ims' { Mime.application_vnd_ms_ims }
        'in' { Mime.text_plain }
        'inc' { Mime.text_x_pascal }
        'ipk' { Mime.application_vnd_shana_informed_package }
        'irm' { Mime.application_vnd_ibm_rights_management }
        'irp' { Mime.application_vnd_irepository_package_xml }
        'iso' { Mime.application_x_iso9660_image }
        'isoimg' { Mime.application_x_iso9660_image }
        'itp' { Mime.application_vnd_shana_informed_formtemplate }
        'ivp' { Mime.application_vnd_immervision_ivp }
        'ivu' { Mime.application_vnd_immervision_ivu }
        'jad' { Mime.text_vnd_sun_j2me_app_descriptor }
        'jam' { Mime.application_vnd_jam }
        'jar' { Mime.application_java_archive }
        'java' { Mime.text_x_java_source }
        'jfi' { Mime.image_pjpeg }
        'jfif' { Mime.image_jpeg }
        'jfif-tbnl' { Mime.image_jpeg }
        'jif' { Mime.image_jpeg }
        'jisp' { Mime.application_vnd_jisp }
        'jlt' { Mime.application_vnd_hp_jlyt }
        'jnlp' { Mime.application_x_java_jnlp_file }
        'joda' { Mime.application_vnd_joost_joda_archive }
        'jpe' { Mime.image_jpeg }
        'jpeg' { Mime.image_jpeg }
        'jpg' { Mime.image_jpeg }
        'jpgm' { Mime.video_jpm }
        'jpgv' { Mime.video_jpeg }
        'jpm' { Mime.video_jpm }
        'js' { Mime.text_javascript }
        'json' { Mime.application_json }
        'k25' { Mime.image_x_kodak_k25 }
        'kar' { Mime.audio_midi }
        'karbon' { Mime.application_vnd_kde_karbon }
        'kdc' { Mime.image_x_kodak_kdc }
        'kfo' { Mime.application_vnd_kde_kformula }
        'kia' { Mime.application_vnd_kidspiration }
        'kil' { Mime.application_x_killustrator }
        'kml' { Mime.application_vnd_google_earth_kml_xml }
        'kmz' { Mime.application_vnd_google_earth_kmz }
        'kne' { Mime.application_vnd_kinar }
        'knp' { Mime.application_vnd_kinar }
        'kon' { Mime.application_vnd_kde_kontour }
        'kpr' { Mime.application_vnd_kde_kpresenter }
        'kpt' { Mime.application_vnd_kde_kpresenter }
        'kra' { Mime.application_x_krita }
        'krz' { Mime.application_x_krita }
        'ksh' { Mime.text_plain }
        'ksp' { Mime.application_vnd_kde_kspread }
        'ktr' { Mime.application_vnd_kahootz }
        'ktz' { Mime.application_vnd_kahootz }
        'kwd' { Mime.application_vnd_kde_kword }
        'kwt' { Mime.application_vnd_kde_kword }
        'latex' { Mime.application_x_latex }
        'lbd' { Mime.application_vnd_llamagraphics_life_balance_desktop }
        'lbe' { Mime.application_vnd_llamagraphics_life_balance_exchange_xml }
        'les' { Mime.application_vnd_hhe_lesson_player }
        'lha' { Mime.application_octet_stream }
        'link66' { Mime.application_vnd_route66_link66_xml }
        'list' { Mime.text_plain }
        'list3820' { Mime.application_vnd_ibm_modcap }
        'listafp' { Mime.application_vnd_ibm_modcap }
        'log' { Mime.text_plain }
        'lostxml' { Mime.application_lost_xml }
        'lrf' { Mime.application_octet_stream }
        'lrm' { Mime.application_vnd_ms_lrm }
        'ltf' { Mime.application_vnd_frogans_ltf }
        'lvp' { Mime.audio_vnd_lucent_voice }
        'lwp' { Mime.application_vnd_lotus_wordpro }
        'lzh' { Mime.application_octet_stream }
        'm13' { Mime.application_x_msmediaview }
        'm14' { Mime.application_x_msmediaview }
        'm1v' { Mime.video_mpeg }
        'm2a' { Mime.audio_mpeg }
        'm2v' { Mime.video_mpeg }
        'm3a' { Mime.audio_mpeg }
        'm3u' { Mime.audio_x_mpegurl }
        'm4a' { Mime.audio_mp4 }
        'm4b' { Mime.audio_mp4 }
        'm4p' { Mime.audio_mp4 }
        'm4r' { Mime.audio_mp4 }
        'm4u' { Mime.video_vnd_mpegurl }
        'm4v' { Mime.audio_mp4 }
        'ma' { Mime.application_mathematica }
        'mag' { Mime.application_vnd_ecowin_chart }
        'maker' { Mime.application_vnd_framemaker }
        'man' { Mime.text_troff }
        'markdn' { Mime.text_markdown }
        'markdown' { Mime.text_markdown }
        'mathml' { Mime.application_mathml_xml }
        'mb' { Mime.application_mathematica }
        'mbk' { Mime.application_vnd_mobius_mbk }
        'mbox' { Mime.application_mbox }
        'mc1' { Mime.application_vnd_medcalcdata }
        'mcd' { Mime.application_vnd_mcd }
        'mcurl' { Mime.text_vnd_curl_mcurl }
        'md' { Mime.text_markdown }
        'mdb' { Mime.application_x_msaccess }
        'mdi' { Mime.image_vnd_ms_modi }
        'mdown' { Mime.text_markdown }
        'me' { Mime.text_troff }
        'mesh' { Mime.model_mesh }
        'mfm' { Mime.application_vnd_mfmp }
        'mgz' { Mime.application_vnd_proteus_magazine }
        'mht' { Mime.message_rfc822 }
        'mhtml' { Mime.message_rfc822 }
        'mid' { Mime.audio_midi }
        'midi' { Mime.audio_midi }
        'mif' { Mime.application_vnd_mif }
        'mime' { Mime.message_rfc822 }
        'mj2' { Mime.video_mj2 }
        'mjp2' { Mime.video_mj2 }
        'mka' { Mime.audio_x_matroska }
        'mkv' { Mime.video_x_matroska }
        'mlp' { Mime.application_vnd_dolby_mlp }
        'mmd' { Mime.application_vnd_chipnuts_karaoke_mmd }
        'mmf' { Mime.application_vnd_smaf }
        'mml' { Mime.application_mathml_xml }
        'mmr' { Mime.image_vnd_fujixerox_edmics_mmr }
        'mny' { Mime.application_x_msmoney }
        'mobi' { Mime.application_x_mobipocket_ebook }
        'mov' { Mime.video_quicktime }
        'movie' { Mime.video_x_sgi_movie }
        'mp2' { Mime.audio_mpeg }
        'mp2a' { Mime.audio_mpeg }
        'mp3' { Mime.audio_mpeg }
        'mp4' { Mime.audio_mp4 }
        'mp4s' { Mime.application_mp4 }
        'mp4v' { Mime.audio_mp4 }
        'mpa' { Mime.video_mpeg }
        'mpc' { Mime.application_vnd_mophun_certificate }
        'mpe' { Mime.video_mpeg }
        'mpeg' { Mime.video_mpeg }
        'mpg' { Mime.video_mpeg }
        'mpg4' { Mime.video_mp4 }
        'mpga' { Mime.audio_mpeg }
        'mpkg' { Mime.application_vnd_apple_installer_xml }
        'mpm' { Mime.application_vnd_blueice_multipass }
        'mpn' { Mime.application_vnd_mophun_application }
        'mpp' { Mime.application_vnd_ms_project }
        'mpt' { Mime.application_vnd_ms_project }
        'mpy' { Mime.application_vnd_ibm_minipay }
        'mqy' { Mime.application_vnd_mobius_mqy }
        'mrc' { Mime.application_marc }
        'mrw' { Mime.image_x_minolta_mrw }
        'ms' { Mime.text_troff }
        'mscml' { Mime.application_mediaservercontrol_xml }
        'mseed' { Mime.application_vnd_fdsn_mseed }
        'mseq' { Mime.application_vnd_mseq }
        'msf' { Mime.application_vnd_epson_msf }
        'msh' { Mime.model_mesh }
        'msi' { Mime.application_x_msdownload }
        'msl' { Mime.application_vnd_mobius_msl }
        'msty' { Mime.application_vnd_muvee_style }
        'mts' { Mime.model_vnd_mts }
        'mus' { Mime.application_vnd_musician }
        'musicxml' { Mime.application_vnd_recordare_musicxml_xml }
        'mvb' { Mime.application_x_msmediaview }
        'mwf' { Mime.application_vnd_mfer }
        'mxf' { Mime.application_mxf }
        'mxl' { Mime.application_vnd_recordare_musicxml }
        'mxml' { Mime.application_xv_xml }
        'mxs' { Mime.application_vnd_triscape_mxs }
        'mxu' { Mime.video_vnd_mpegurl }
        'n-gage' { Mime.application_vnd_nokia_n_gage_symbian_install }
        'nb' { Mime.application_mathematica }
        'nc' { Mime.application_x_netcdf }
        'ncx' { Mime.application_x_dtbncx_xml }
        'nef' { Mime.image_x_nikon_nef }
        'ngdat' { Mime.application_vnd_nokia_n_gage_data }
        'nlu' { Mime.application_vnd_neurolanguage_nlu }
        'nml' { Mime.application_vnd_enliven }
        'nnd' { Mime.application_vnd_noblenet_directory }
        'nns' { Mime.application_vnd_noblenet_sealer }
        'nnw' { Mime.application_vnd_noblenet_web }
        'npx' { Mime.image_vnd_net_fpx }
        'nsf' { Mime.application_vnd_lotus_notes }
        'nws' { Mime.message_rfc822 }
        'o' { Mime.application_octet_stream }
        'oa2' { Mime.application_vnd_fujitsu_oasys2 }
        'oa3' { Mime.application_vnd_fujitsu_oasys3 }
        'oas' { Mime.application_vnd_fujitsu_oasys }
        'obd' { Mime.application_x_msbinder }
        'obj' { Mime.application_octet_stream }
        'oda' { Mime.application_oda }
        'odb' { Mime.application_vnd_oasis_opendocument_database }
        'odc' { Mime.application_vnd_oasis_opendocument_chart }
        'odf' { Mime.application_vnd_oasis_opendocument_formula }
        'odft' { Mime.application_vnd_oasis_opendocument_formula_template }
        'odg' { Mime.application_vnd_oasis_opendocument_graphics }
        'odi' { Mime.application_vnd_oasis_opendocument_image }
        'odp' { Mime.application_vnd_oasis_opendocument_presentation }
        'ods' { Mime.application_vnd_oasis_opendocument_spreadsheet }
        'odt' { Mime.application_vnd_oasis_opendocument_text }
        'oga' { Mime.audio_ogg }
        'ogg' { Mime.audio_ogg }
        'ogv' { Mime.video_ogg }
        'ogx' { Mime.application_ogg }
        'onepkg' { Mime.application_onenote }
        'onetmp' { Mime.application_onenote }
        'onetoc' { Mime.application_onenote }
        'onetoc2' { Mime.application_onenote }
        'opf' { Mime.application_oebps_package_xml }
        'oprc' { Mime.application_vnd_palm }
        'opus' { Mime.audio_opus }
        'orf' { Mime.image_x_olympus_orf }
        'org' { Mime.application_vnd_lotus_organizer }
        'osf' { Mime.application_vnd_yamaha_openscoreformat }
        'osfpvg' { Mime.application_vnd_yamaha_openscoreformat_osfpvg_xml }
        'otc' { Mime.application_vnd_oasis_opendocument_chart_template }
        'otf' { Mime.application_x_font_otf }
        'otg' { Mime.application_vnd_oasis_opendocument_graphics_template }
        'oth' { Mime.application_vnd_oasis_opendocument_text_web }
        'oti' { Mime.application_vnd_oasis_opendocument_image_template }
        'otm' { Mime.application_vnd_oasis_opendocument_text_master }
        'otp' { Mime.application_vnd_oasis_opendocument_presentation_template }
        'ots' { Mime.application_vnd_oasis_opendocument_spreadsheet_template }
        'ott' { Mime.application_vnd_oasis_opendocument_text_template }
        'oxt' { Mime.application_vnd_openofficeorg_extension }
        'p' { Mime.text_x_pascal }
        'p10' { Mime.application_pkcs10 }
        'p12' { Mime.application_x_pkcs12 }
        'p7b' { Mime.application_x_pkcs7_certificates }
        'p7c' { Mime.application_pkcs7_mime }
        'p7m' { Mime.application_pkcs7_mime }
        'p7r' { Mime.application_x_pkcs7_certreqresp }
        'p7s' { Mime.application_pkcs7_signature }
        'pas' { Mime.text_x_pascal }
        'pbd' { Mime.application_vnd_powerbuilder6 }
        'pbm' { Mime.image_x_portable_bitmap }
        'pcf' { Mime.application_x_font_pcf }
        'pcl' { Mime.application_vnd_hp_pcl }
        'pclxl' { Mime.application_vnd_hp_pclxl }
        'pct' { Mime.image_x_pict }
        'pcurl' { Mime.application_vnd_curl_pcurl }
        'pcx' { Mime.image_x_pcx }
        'pdb' { Mime.application_vnd_palm }
        'pdf' { Mime.application_pdf }
        'pef' { Mime.image_x_pentax_pef }
        'pfa' { Mime.application_x_font_type1 }
        'pfb' { Mime.application_x_font_type1 }
        'pfm' { Mime.application_x_font_type1 }
        'pfr' { Mime.application_font_tdpfr }
        'pfx' { Mime.application_x_pkcs12 }
        'pgm' { Mime.image_x_portable_graymap }
        'pgn' { Mime.application_x_chess_pgn }
        'pgp' { Mime.application_pgp_encrypted }
        'pic' { Mime.image_x_pict }
        'pjpg' { Mime.image_jpeg }
        'pkg' { Mime.application_octet_stream }
        'pki' { Mime.application_pkixcmp }
        'pkipath' { Mime.application_pkix_pkipath }
        'pl' { Mime.text_plain }
        'plb' { Mime.application_vnd_3gpp_pic_bw_large }
        'plc' { Mime.application_vnd_mobius_plc }
        'plf' { Mime.application_vnd_pocketlearn }
        'pls' { Mime.application_pls_xml }
        'pm' { Mime.application_x_perl }
        'pml' { Mime.application_vnd_ctc_posml }
        'png' { Mime.image_png }
        'pnm' { Mime.image_x_portable_anymap }
        'portpkg' { Mime.application_vnd_macports_portpkg }
        'pot' { Mime.application_vnd_ms_powerpoint }
        'potm' { Mime.application_vnd_ms_powerpoint_template_macroenabled_12 }
        'potx' { Mime.application_vnd_openxmlformats_officedocument_presentationml_template }
        'pp' { Mime.text_x_pascal }
        'ppa' { Mime.application_vnd_ms_powerpoint }
        'ppam' { Mime.application_vnd_ms_powerpoint_addin_macroenabled_12 }
        'ppd' { Mime.application_vnd_cups_ppd }
        'ppm' { Mime.image_x_portable_pixmap }
        'pps' { Mime.application_vnd_ms_powerpoint }
        'ppsm' { Mime.application_vnd_ms_powerpoint_slideshow_macroenabled_12 }
        'ppsx' { Mime.application_vnd_openxmlformats_officedocument_presentationml_slideshow }
        'ppt' { Mime.application_vnd_ms_powerpoint }
        'pptm' { Mime.application_vnd_ms_powerpoint_presentation_macroenabled_12 }
        'pptx' { Mime.application_vnd_openxmlformats_officedocument_presentationml_presentation }
        'pqa' { Mime.application_vnd_palm }
        'prc' { Mime.application_x_mobipocket_ebook }
        'pre' { Mime.application_vnd_lotus_freelance }
        'prf' { Mime.application_pics_rules }
        'prql' { Mime.application_prql }
        'ps' { Mime.application_postscript }
        'psb' { Mime.application_vnd_3gpp_pic_bw_small }
        'psd' { Mime.image_vnd_adobe_photoshop }
        'psf' { Mime.application_x_font_linux_psf }
        'ptid' { Mime.application_vnd_pvi_ptid1 }
        'ptx' { Mime.image_x_pentax_pef }
        'pub' { Mime.application_x_mspublisher }
        'pvb' { Mime.application_vnd_3gpp_pic_bw_var }
        'pwn' { Mime.application_vnd_3m_post_it_notes }
        'pwz' { Mime.application_vnd_ms_powerpoint }
        'py' { Mime.text_x_python }
        'pya' { Mime.audio_vnd_ms_playready_media_pya }
        'pyc' { Mime.text_x_python }
        'pyd' { Mime.text_x_python }
        'pyo' { Mime.text_x_python }
        'pyv' { Mime.video_vnd_ms_playready_media_pyv }
        'qam' { Mime.application_vnd_epson_quickanime }
        'qbo' { Mime.application_vnd_intu_qbo }
        'qfx' { Mime.application_vnd_intu_qfx }
        'qps' { Mime.application_vnd_publishare_delta_tree }
        'qt' { Mime.video_quicktime }
        'qwd' { Mime.application_vnd_quark_quarkxpress }
        'qwt' { Mime.application_vnd_quark_quarkxpress }
        'qxb' { Mime.application_vnd_quark_quarkxpress }
        'qxd' { Mime.application_vnd_quark_quarkxpress }
        'qxl' { Mime.application_vnd_quark_quarkxpress }
        'qxt' { Mime.application_vnd_quark_quarkxpress }
        'ra' { Mime.audio_x_pn_realaudio }
        'raf' { Mime.image_x_fuji_raf }
        'ram' { Mime.audio_x_pn_realaudio }
        'rar' { Mime.application_vnd_rar }
        'ras' { Mime.image_x_cmu_raster }
        'raw' { Mime.image_x_panasonic_raw }
        'rcprofile' { Mime.application_vnd_ipunplugged_rcprofile }
        'rdf' { Mime.application_rdf_xml }
        'rdz' { Mime.application_vnd_data_vision_rdz }
        'rep' { Mime.application_vnd_businessobjects }
        'res' { Mime.application_x_dtbresource_xml }
        'rgb' { Mime.image_x_rgb }
        'rif' { Mime.application_reginfo_xml }
        'rl' { Mime.application_resource_lists_xml }
        'rlc' { Mime.image_vnd_fujixerox_edmics_rlc }
        'rld' { Mime.application_resource_lists_diff_xml }
        'rm' { Mime.application_vnd_rn_realmedia }
        'rmi' { Mime.audio_midi }
        'rmp' { Mime.audio_x_pn_realaudio_plugin }
        'rms' { Mime.application_vnd_jcp_javame_midlet_rms }
        'rnc' { Mime.application_relax_ng_compact_syntax }
        'roff' { Mime.text_troff }
        'rpa' { Mime.application_x_redhat_package_manager }
        'rpm' { Mime.application_x_rpm }
        'rpss' { Mime.application_vnd_nokia_radio_presets }
        'rpst' { Mime.application_vnd_nokia_radio_preset }
        'rq' { Mime.application_sparql_query }
        'rs' { Mime.application_rls_services_xml }
        'rsd' { Mime.application_rsd_xml }
        'rss' { Mime.application_rss_xml }
        'rtf' { Mime.application_rtf }
        'rtx' { Mime.text_richtext }
        'rw2' { Mime.image_x_panasonic_raw }
        'rwl' { Mime.image_x_panasonic_raw }
        's' { Mime.text_x_asm }
        'saf' { Mime.application_vnd_yamaha_smaf_audio }
        'sbml' { Mime.application_sbml_xml }
        'sc' { Mime.application_vnd_ibm_secure_container }
        'scd' { Mime.application_x_msschedule }
        'scm' { Mime.application_vnd_lotus_screencam }
        'scq' { Mime.application_scvp_cv_request }
        'scs' { Mime.application_scvp_cv_response }
        'scurl' { Mime.text_vnd_curl_scurl }
        'sda' { Mime.application_vnd_stardivision_draw }
        'sdc' { Mime.application_vnd_stardivision_calc }
        'sdd' { Mime.application_vnd_stardivision_impress }
        'sdkd' { Mime.application_vnd_solent_sdkm_xml }
        'sdkm' { Mime.application_vnd_solent_sdkm_xml }
        'sdp' { Mime.application_sdp }
        'sdw' { Mime.application_vnd_stardivision_writer }
        'see' { Mime.application_vnd_seemail }
        'seed' { Mime.application_vnd_fdsn_seed }
        'sema' { Mime.application_vnd_sema }
        'semd' { Mime.application_vnd_semd }
        'semf' { Mime.application_vnd_semf }
        'ser' { Mime.application_java_serialized_object }
        'setpay' { Mime.application_set_payment_initiation }
        'setreg' { Mime.application_set_registration_initiation }
        'sfd-hdstx' { Mime.application_vnd_hydrostatix_sof_data }
        'sfs' { Mime.application_vnd_spotfire_sfs }
        'sgl' { Mime.application_vnd_stardivision_writer_global }
        'sgm' { Mime.text_sgml }
        'sgml' { Mime.text_sgml }
        'sh' { Mime.application_x_shellscript }
        'shar' { Mime.application_x_shar }
        'shf' { Mime.application_shf_xml }
        'si' { Mime.text_vnd_wap_si }
        'sic' { Mime.application_vnd_wap_sic }
        'sig' { Mime.application_pgp_signature }
        'silo' { Mime.model_mesh }
        'sis' { Mime.application_vnd_symbian_install }
        'sisx' { Mime.application_vnd_symbian_install }
        'sit' { Mime.application_x_stuffit }
        'sitx' { Mime.application_x_stuffitx }
        'skd' { Mime.application_vnd_koan }
        'skm' { Mime.application_vnd_koan }
        'skp' { Mime.application_vnd_koan }
        'skt' { Mime.application_vnd_koan }
        'sl' { Mime.text_vnd_wap_sl }
        'slc' { Mime.application_vnd_wap_slc }
        'sldm' { Mime.application_vnd_ms_powerpoint_slide_macroenabled_12 }
        'sldx' { Mime.application_vnd_openxmlformats_officedocument_presentationml_slide }
        'slt' { Mime.application_vnd_epson_salt }
        'smf' { Mime.application_vnd_stardivision_math }
        'smi' { Mime.application_smil_xml }
        'smil' { Mime.application_smil_xml }
        'snd' { Mime.audio_basic }
        'snf' { Mime.application_x_font_snf }
        'so' { Mime.application_octet_stream }
        'spc' { Mime.application_x_pkcs7_certificates }
        'spf' { Mime.application_vnd_yamaha_smaf_phrase }
        'spl' { Mime.application_x_futuresplash }
        'spot' { Mime.text_vnd_in3d_spot }
        'spp' { Mime.application_scvp_vp_response }
        'spq' { Mime.application_scvp_vp_request }
        'spx' { Mime.audio_ogg }
        'sqlite' { Mime.application_vnd_sqlite3 }
        'sqlite-shm' { Mime.application_vnd_sqlite3 }
        'sqlite-wal' { Mime.application_vnd_sqlite3 }
        'sqlite3' { Mime.application_vnd_sqlite3 }
        'sr2' { Mime.image_x_sony_sr2 }
        'src' { Mime.application_x_wais_source }
        'srf' { Mime.image_x_sony_srf }
        'srx' { Mime.application_sparql_results_xml }
        'sse' { Mime.application_vnd_kodak_descriptor }
        'ssf' { Mime.application_vnd_epson_ssf }
        'ssml' { Mime.application_ssml_xml }
        'stc' { Mime.application_vnd_sun_xml_calc_template }
        'std' { Mime.application_vnd_sun_xml_draw_template }
        'stf' { Mime.application_vnd_wt_stf }
        'sti' { Mime.application_vnd_sun_xml_impress_template }
        'stk' { Mime.application_hyperstudio }
        'stl' { Mime.application_vnd_ms_pki_stl }
        'str' { Mime.application_vnd_pg_format }
        'stw' { Mime.application_vnd_sun_xml_writer_template }
        'sus' { Mime.application_vnd_sus_calendar }
        'susp' { Mime.application_vnd_sus_calendar }
        'sv4cpio' { Mime.application_x_sv4cpio }
        'sv4crc' { Mime.application_x_sv4crc }
        'svd' { Mime.application_vnd_svd }
        'svg' { Mime.image_svg_xml }
        'svgz' { Mime.image_svg_xml }
        'swa' { Mime.application_x_director }
        'swf' { Mime.application_x_shockwave_flash }
        'swi' { Mime.application_vnd_arastra_swi }
        'sxc' { Mime.application_vnd_sun_xml_calc }
        'sxd' { Mime.application_vnd_sun_xml_draw }
        'sxg' { Mime.application_vnd_sun_xml_writer_global }
        'sxi' { Mime.application_vnd_sun_xml_impress }
        'sxm' { Mime.application_vnd_sun_xml_math }
        'sxw' { Mime.application_vnd_sun_xml_writer }
        't' { Mime.text_troff }
        'tao' { Mime.application_vnd_tao_intent_module_archive }
        'tar' { Mime.application_x_tar }
        'tcap' { Mime.application_vnd_3gpp2_tcap }
        'tcl' { Mime.application_x_tcl }
        'teacher' { Mime.application_vnd_smart_teacher }
        'test' { Mime.test_mimetype }
        'tex' { Mime.application_x_tex }
        'texi' { Mime.application_x_texinfo }
        'texinfo' { Mime.application_x_texinfo }
        'text' { Mime.text_plain }
        'tfm' { Mime.application_x_tex_tfm }
        'tgz' { Mime.application_x_gzip }
        'tif' { Mime.image_tiff }
        'tiff' { Mime.image_tiff }
        'tmo' { Mime.application_vnd_tmobile_livetv }
        'torrent' { Mime.application_x_bittorrent }
        'tpl' { Mime.application_vnd_groove_tool_template }
        'tpt' { Mime.application_vnd_trid_tpt }
        'tr' { Mime.text_troff }
        'tra' { Mime.application_vnd_trueapp }
        'trm' { Mime.application_x_msterminal }
        'ts' { Mime.video_mp2t }
        'tsv' { Mime.text_tab_separated_values }
        'ttc' { Mime.application_x_font_ttf }
        'ttf' { Mime.application_x_font_ttf }
        'twd' { Mime.application_vnd_simtech_mindmapper }
        'twds' { Mime.application_vnd_simtech_mindmapper }
        'txd' { Mime.application_vnd_genomatix_tuxedo }
        'txf' { Mime.application_vnd_mobius_txf }
        'txt' { Mime.text_plain }
        'u32' { Mime.application_x_authorware_bin }
        'udeb' { Mime.application_vnd_debian_binary_package }
        'ufd' { Mime.application_vnd_ufdl }
        'ufdl' { Mime.application_vnd_ufdl }
        'umj' { Mime.application_vnd_umajin }
        'unityweb' { Mime.application_vnd_unity }
        'uoml' { Mime.application_vnd_uoml_xml }
        'uri' { Mime.text_uri_list }
        'uris' { Mime.text_uri_list }
        'urls' { Mime.text_uri_list }
        'ustar' { Mime.application_x_ustar }
        'utz' { Mime.application_vnd_uiq_theme }
        'uu' { Mime.text_x_uuencode }
        'vcd' { Mime.application_x_cdlink }
        'vcf' { Mime.text_x_vcard }
        'vcg' { Mime.application_vnd_groove_vcard }
        'vcs' { Mime.text_x_vcalendar }
        'vcx' { Mime.application_vnd_vcx }
        'vis' { Mime.application_vnd_visionary }
        'viv' { Mime.video_vnd_vivo }
        'vor' { Mime.application_vnd_stardivision_writer }
        'vox' { Mime.application_x_authorware_bin }
        'vrml' { Mime.model_vrml }
        'vsd' { Mime.application_vnd_visio }
        'vsdx' { Mime.application_vnd_visio }
        'vsf' { Mime.application_vnd_vsf }
        'vss' { Mime.application_vnd_visio }
        'vssm' { Mime.application_vnd_visio }
        'vssx' { Mime.application_vnd_visio }
        'vst' { Mime.application_vnd_visio }
        'vstm' { Mime.application_vnd_visio }
        'vstx' { Mime.application_vnd_visio }
        'vsw' { Mime.application_vnd_visio }
        'vtu' { Mime.model_vnd_vtu }
        'vxml' { Mime.application_voicexml_xml }
        'w3d' { Mime.application_x_director }
        'wad' { Mime.application_x_doom }
        'wasm' { Mime.application_wasm }
        'wav' { Mime.audio_vnd_wav }
        'wax' { Mime.audio_x_ms_wax }
        'wbmp' { Mime.image_vnd_wap_wbmp }
        'wbs' { Mime.application_vnd_criticaltools_wbs_xml }
        'wbxml' { Mime.application_vnd_wap_wbxml }
        'wcm' { Mime.application_vnd_ms_works }
        'wdb' { Mime.application_vnd_ms_works }
        'weba' { Mime.audio_webm }
        'webm' { Mime.video_webm }
        'webp' { Mime.image_webp }
        'whl' { Mime.text_x_python }
        'wiz' { Mime.application_msword }
        'wks' { Mime.application_vnd_ms_works }
        'wm' { Mime.video_x_ms_wm }
        'wma' { Mime.audio_x_ms_wma }
        'wmd' { Mime.application_x_ms_wmd }
        'wmf' { Mime.application_x_msmetafile }
        'wml' { Mime.text_vnd_wap_wml }
        'wmlc' { Mime.application_vnd_wap_wmlc }
        'wmls' { Mime.text_vnd_wap_wmlscript }
        'wmlsc' { Mime.application_vnd_wap_wmlscriptc }
        'wmv' { Mime.video_x_ms_wmv }
        'wmx' { Mime.video_x_ms_wmx }
        'wmz' { Mime.application_x_ms_wmz }
        'woff' { Mime.font_woff }
        'woff2' { Mime.font_woff2 }
        'wpd' { Mime.application_vnd_wordperfect }
        'wpl' { Mime.application_vnd_ms_wpl }
        'wps' { Mime.application_vnd_ms_works }
        'wqd' { Mime.application_vnd_wqd }
        'wri' { Mime.application_x_mswrite }
        'wrl' { Mime.model_vrml }
        'wsdl' { Mime.application_wsdl_xml }
        'wspolicy' { Mime.application_wspolicy_xml }
        'wtb' { Mime.application_vnd_webturbo }
        'wvx' { Mime.video_x_ms_wvx }
        'x32' { Mime.application_x_authorware_bin }
        'x3d' { Mime.application_vnd_hzn_3d_crossword }
        'x3f' { Mime.image_x_sigma_x3f }
        'xap' { Mime.application_x_silverlight_app }
        'xar' { Mime.application_vnd_xara }
        'xbap' { Mime.application_x_ms_xbap }
        'xbd' { Mime.application_vnd_fujixerox_docuworks_binder }
        'xbm' { Mime.image_x_xbitmap }
        'xdm' { Mime.application_vnd_syncml_dm_xml }
        'xdp' { Mime.application_vnd_adobe_xdp_xml }
        'xdw' { Mime.application_vnd_fujixerox_docuworks }
        'xenc' { Mime.application_xenc_xml }
        'xer' { Mime.application_patch_ops_error_xml }
        'xfdf' { Mime.application_vnd_adobe_xfdf }
        'xfdl' { Mime.application_vnd_xfdl }
        'xht' { Mime.application_xhtml_xml }
        'xhtml' { Mime.application_xhtml_xml }
        'xhvml' { Mime.application_xv_xml }
        'xif' { Mime.image_vnd_xiff }
        'xla' { Mime.application_vnd_ms_excel }
        'xlam' { Mime.application_vnd_ms_excel_addin_macroenabled_12 }
        'xlb' { Mime.application_vnd_ms_excel }
        'xlc' { Mime.application_vnd_ms_excel }
        'xlm' { Mime.application_vnd_ms_excel }
        'xls' { Mime.application_vnd_ms_excel }
        'xlsb' { Mime.application_vnd_ms_excel_sheet_binary_macroenabled_12 }
        'xlsm' { Mime.application_vnd_ms_excel_sheet_macroenabled_12 }
        'xlsx' { Mime.application_vnd_openxmlformats_officedocument_spreadsheetml_sheet }
        'xlt' { Mime.application_vnd_ms_excel }
        'xltm' { Mime.application_vnd_ms_excel_template_macroenabled_12 }
        'xltx' { Mime.application_vnd_openxmlformats_officedocument_spreadsheetml_template }
        'xlw' { Mime.application_vnd_ms_excel }
        'xml' { Mime.application_rss_xml }
        'xo' { Mime.application_vnd_olpc_sugar }
        'xop' { Mime.application_xop_xml }
        'xpdl' { Mime.application_xml }
        'xpi' { Mime.application_x_xpinstall }
        'xpm' { Mime.image_x_xpixmap }
        'xpr' { Mime.application_vnd_is_xpr }
        'xps' { Mime.application_vnd_ms_xpsdocument }
        'xpw' { Mime.application_vnd_intercon_formnet }
        'xpx' { Mime.application_vnd_intercon_formnet }
        'xsl' { Mime.application_xml }
        'xslt' { Mime.application_xslt_xml }
        'xsm' { Mime.application_vnd_syncml_xml }
        'xspf' { Mime.application_xspf_xml }
        'xul' { Mime.application_vnd_mozilla_xul_xml }
        'xvm' { Mime.application_xv_xml }
        'xvml' { Mime.application_xv_xml }
        'xwd' { Mime.image_x_xwindowdump }
        'xyz' { Mime.chemical_x_xyz }
        'yaml' { Mime.application_yaml }
        'yml' { Mime.application_yaml }
        'zabw' { Mime.application_x_abiword }
        'zaz' { Mime.application_vnd_zzazz_deck_xml }
        'zip' { Mime.application_zip }
        'zir' { Mime.application_vnd_zul }
        'zirz' { Mime.application_vnd_zul }
        'zmm' { Mime.application_vnd_handheld_entertainment_xml }
        else { none }
    }
}
