module mime

/*
https://www.iana.org/assignments/media-types/media-types.xhtml
*/
pub enum Mime {
	application_javascript
	application_json
	image_avif
	image_jpeg
	image_png
	image_webp
	svg_xml
	text_css
	text_html
}
